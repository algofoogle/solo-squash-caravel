magic
tech sky130A
magscale 1 2
timestamp 1679986742
<< viali >>
rect 7205 37281 7239 37315
rect 1777 37213 1811 37247
rect 7481 37213 7515 37247
rect 14289 37213 14323 37247
rect 20269 37213 20303 37247
rect 27169 37213 27203 37247
rect 32965 37213 32999 37247
rect 38025 37213 38059 37247
rect 1593 37077 1627 37111
rect 14473 37077 14507 37111
rect 20085 37077 20119 37111
rect 27353 37077 27387 37111
rect 33149 37077 33183 37111
rect 38209 37077 38243 37111
rect 19441 36873 19475 36907
rect 19625 36737 19659 36771
rect 1593 34561 1627 34595
rect 1777 34357 1811 34391
rect 14657 34017 14691 34051
rect 9873 33949 9907 33983
rect 12357 33949 12391 33983
rect 13737 33949 13771 33983
rect 14381 33949 14415 33983
rect 14473 33949 14507 33983
rect 15945 33949 15979 33983
rect 16129 33949 16163 33983
rect 12541 33881 12575 33915
rect 9689 33813 9723 33847
rect 13553 33813 13587 33847
rect 14657 33813 14691 33847
rect 16037 33813 16071 33847
rect 16129 33609 16163 33643
rect 9842 33541 9876 33575
rect 7748 33473 7782 33507
rect 12633 33473 12667 33507
rect 14269 33473 14303 33507
rect 15853 33473 15887 33507
rect 7481 33405 7515 33439
rect 9597 33405 9631 33439
rect 12357 33405 12391 33439
rect 14013 33405 14047 33439
rect 16129 33405 16163 33439
rect 15393 33337 15427 33371
rect 8861 33269 8895 33303
rect 10977 33269 11011 33303
rect 15945 33269 15979 33303
rect 8585 33065 8619 33099
rect 7297 32929 7331 32963
rect 8217 32929 8251 32963
rect 9137 32929 9171 32963
rect 15577 32929 15611 32963
rect 16037 32929 16071 32963
rect 7481 32861 7515 32895
rect 8401 32861 8435 32895
rect 9413 32861 9447 32895
rect 10885 32861 10919 32895
rect 11161 32861 11195 32895
rect 12173 32861 12207 32895
rect 14749 32861 14783 32895
rect 14841 32861 14875 32895
rect 16293 32861 16327 32895
rect 38301 32861 38335 32895
rect 12440 32793 12474 32827
rect 14565 32793 14599 32827
rect 15393 32793 15427 32827
rect 7665 32725 7699 32759
rect 13553 32725 13587 32759
rect 14841 32725 14875 32759
rect 17417 32725 17451 32759
rect 8401 32521 8435 32555
rect 12725 32521 12759 32555
rect 13645 32521 13679 32555
rect 17233 32521 17267 32555
rect 13461 32453 13495 32487
rect 6561 32385 6595 32419
rect 6828 32385 6862 32419
rect 8585 32385 8619 32419
rect 9413 32385 9447 32419
rect 10241 32385 10275 32419
rect 10425 32385 10459 32419
rect 10885 32385 10919 32419
rect 11069 32385 11103 32419
rect 11897 32385 11931 32419
rect 12909 32385 12943 32419
rect 13737 32385 13771 32419
rect 15669 32385 15703 32419
rect 15853 32385 15887 32419
rect 15945 32385 15979 32419
rect 17049 32385 17083 32419
rect 17877 32385 17911 32419
rect 9321 32317 9355 32351
rect 11805 32317 11839 32351
rect 14197 32317 14231 32351
rect 15761 32317 15795 32351
rect 16865 32317 16899 32351
rect 9781 32249 9815 32283
rect 13461 32249 13495 32283
rect 7941 32181 7975 32215
rect 10333 32181 10367 32215
rect 10977 32181 11011 32215
rect 12173 32181 12207 32215
rect 14427 32181 14461 32215
rect 15485 32181 15519 32215
rect 17693 32181 17727 32215
rect 8401 31977 8435 32011
rect 9505 31977 9539 32011
rect 13001 31977 13035 32011
rect 13185 31977 13219 32011
rect 14841 31977 14875 32011
rect 5181 31909 5215 31943
rect 8585 31909 8619 31943
rect 18061 31909 18095 31943
rect 9873 31841 9907 31875
rect 10333 31841 10367 31875
rect 11897 31841 11931 31875
rect 15485 31841 15519 31875
rect 15578 31841 15612 31875
rect 15669 31841 15703 31875
rect 16681 31841 16715 31875
rect 2605 31773 2639 31807
rect 2881 31773 2915 31807
rect 5181 31773 5215 31807
rect 5365 31773 5399 31807
rect 5825 31773 5859 31807
rect 6009 31773 6043 31807
rect 6469 31773 6503 31807
rect 6745 31773 6779 31807
rect 9413 31773 9447 31807
rect 10609 31773 10643 31807
rect 10885 31773 10919 31807
rect 11529 31773 11563 31807
rect 11621 31773 11655 31807
rect 14289 31773 14323 31807
rect 14657 31773 14691 31807
rect 15761 31773 15795 31807
rect 16948 31773 16982 31807
rect 19993 31773 20027 31807
rect 8217 31705 8251 31739
rect 8417 31705 8451 31739
rect 11989 31705 12023 31739
rect 12817 31705 12851 31739
rect 14473 31705 14507 31739
rect 14565 31705 14599 31739
rect 5917 31637 5951 31671
rect 10517 31637 10551 31671
rect 10701 31637 10735 31671
rect 11345 31637 11379 31671
rect 13017 31637 13051 31671
rect 15301 31637 15335 31671
rect 19809 31637 19843 31671
rect 6745 31433 6779 31467
rect 10517 31433 10551 31467
rect 12449 31433 12483 31467
rect 22477 31433 22511 31467
rect 23305 31433 23339 31467
rect 10793 31365 10827 31399
rect 11003 31365 11037 31399
rect 13277 31365 13311 31399
rect 20076 31365 20110 31399
rect 24409 31365 24443 31399
rect 3801 31297 3835 31331
rect 4077 31297 4111 31331
rect 5273 31297 5307 31331
rect 6653 31297 6687 31331
rect 6837 31297 6871 31331
rect 7297 31297 7331 31331
rect 7481 31297 7515 31331
rect 8171 31297 8205 31331
rect 8306 31297 8340 31331
rect 8406 31297 8440 31331
rect 8585 31297 8619 31331
rect 9597 31297 9631 31331
rect 9689 31297 9723 31331
rect 9873 31297 9907 31331
rect 10701 31297 10735 31331
rect 10885 31297 10919 31331
rect 11897 31297 11931 31331
rect 12265 31297 12299 31331
rect 13093 31297 13127 31331
rect 13185 31297 13219 31331
rect 15117 31297 15151 31331
rect 16313 31297 16347 31331
rect 17325 31297 17359 31331
rect 18225 31297 18259 31331
rect 22017 31297 22051 31331
rect 23121 31297 23155 31331
rect 23397 31297 23431 31331
rect 2513 31229 2547 31263
rect 2789 31229 2823 31263
rect 5365 31229 5399 31263
rect 9965 31229 9999 31263
rect 11161 31229 11195 31263
rect 11805 31229 11839 31263
rect 13461 31229 13495 31263
rect 14841 31229 14875 31263
rect 17969 31229 18003 31263
rect 19809 31229 19843 31263
rect 24593 31229 24627 31263
rect 24777 31229 24811 31263
rect 12909 31161 12943 31195
rect 17509 31161 17543 31195
rect 24409 31161 24443 31195
rect 5641 31093 5675 31127
rect 7297 31093 7331 31127
rect 7941 31093 7975 31127
rect 10057 31093 10091 31127
rect 12173 31093 12207 31127
rect 16129 31093 16163 31127
rect 19349 31093 19383 31127
rect 21189 31093 21223 31127
rect 22293 31093 22327 31127
rect 22937 31093 22971 31127
rect 24685 31093 24719 31127
rect 11897 30889 11931 30923
rect 12541 30889 12575 30923
rect 14657 30889 14691 30923
rect 15485 30889 15519 30923
rect 15669 30889 15703 30923
rect 16313 30889 16347 30923
rect 16497 30889 16531 30923
rect 17877 30889 17911 30923
rect 18705 30889 18739 30923
rect 19809 30889 19843 30923
rect 24593 30889 24627 30923
rect 6561 30821 6595 30855
rect 18889 30821 18923 30855
rect 23489 30821 23523 30855
rect 24961 30821 24995 30855
rect 2421 30753 2455 30787
rect 5917 30753 5951 30787
rect 6101 30753 6135 30787
rect 10609 30753 10643 30787
rect 11437 30753 11471 30787
rect 12725 30753 12759 30787
rect 17233 30753 17267 30787
rect 20913 30753 20947 30787
rect 21189 30753 21223 30787
rect 23029 30753 23063 30787
rect 2697 30685 2731 30719
rect 4629 30685 4663 30719
rect 4813 30685 4847 30719
rect 4905 30685 4939 30719
rect 5825 30685 5859 30719
rect 6837 30685 6871 30719
rect 7757 30685 7791 30719
rect 7849 30685 7883 30719
rect 8033 30685 8067 30719
rect 8125 30685 8159 30719
rect 9413 30685 9447 30719
rect 9597 30685 9631 30719
rect 9689 30685 9723 30719
rect 10205 30685 10239 30719
rect 10333 30685 10367 30719
rect 10425 30679 10459 30713
rect 11161 30685 11195 30719
rect 11345 30685 11379 30719
rect 11529 30685 11563 30719
rect 11713 30685 11747 30719
rect 12817 30685 12851 30719
rect 13185 30685 13219 30719
rect 17049 30685 17083 30719
rect 18061 30685 18095 30719
rect 20453 30685 20487 30719
rect 23121 30685 23155 30719
rect 24777 30685 24811 30719
rect 25053 30685 25087 30719
rect 16359 30651 16393 30685
rect 6101 30617 6135 30651
rect 6561 30617 6595 30651
rect 9229 30617 9263 30651
rect 14473 30617 14507 30651
rect 15301 30617 15335 30651
rect 15511 30617 15545 30651
rect 16129 30617 16163 30651
rect 18521 30617 18555 30651
rect 19441 30617 19475 30651
rect 19625 30617 19659 30651
rect 4445 30549 4479 30583
rect 6745 30549 6779 30583
rect 7573 30549 7607 30583
rect 12863 30549 12897 30583
rect 13093 30549 13127 30583
rect 14673 30549 14707 30583
rect 14841 30549 14875 30583
rect 18721 30549 18755 30583
rect 20269 30549 20303 30583
rect 3801 30345 3835 30379
rect 4445 30345 4479 30379
rect 5825 30345 5859 30379
rect 8493 30345 8527 30379
rect 9689 30345 9723 30379
rect 10517 30345 10551 30379
rect 12909 30345 12943 30379
rect 16313 30345 16347 30379
rect 18981 30345 19015 30379
rect 22477 30345 22511 30379
rect 23765 30345 23799 30379
rect 6837 30277 6871 30311
rect 7573 30277 7607 30311
rect 12633 30277 12667 30311
rect 14197 30277 14231 30311
rect 14565 30277 14599 30311
rect 16129 30277 16163 30311
rect 22017 30277 22051 30311
rect 25329 30277 25363 30311
rect 2688 30209 2722 30243
rect 4386 30209 4420 30243
rect 5549 30209 5583 30243
rect 6561 30209 6595 30243
rect 6653 30209 6687 30243
rect 7481 30209 7515 30243
rect 8309 30209 8343 30243
rect 9229 30209 9263 30243
rect 10333 30209 10367 30243
rect 10517 30209 10551 30243
rect 10977 30209 11011 30243
rect 12750 30209 12784 30243
rect 13553 30209 13587 30243
rect 14381 30209 14415 30243
rect 14473 30209 14507 30243
rect 15761 30209 15795 30243
rect 16865 30209 16899 30243
rect 17121 30209 17155 30243
rect 18889 30209 18923 30243
rect 19073 30209 19107 30243
rect 20085 30209 20119 30243
rect 20352 30209 20386 30243
rect 23397 30209 23431 30243
rect 2421 30141 2455 30175
rect 4905 30141 4939 30175
rect 5825 30141 5859 30175
rect 6837 30141 6871 30175
rect 8125 30141 8159 30175
rect 12265 30141 12299 30175
rect 12541 30141 12575 30175
rect 13737 30141 13771 30175
rect 23305 30141 23339 30175
rect 24685 30141 24719 30175
rect 25053 30141 25087 30175
rect 25145 30141 25179 30175
rect 5641 30073 5675 30107
rect 22293 30073 22327 30107
rect 4261 30005 4295 30039
rect 4813 30005 4847 30039
rect 9321 30005 9355 30039
rect 11069 30005 11103 30039
rect 14749 30005 14783 30039
rect 16129 30005 16163 30039
rect 18245 30005 18279 30039
rect 21465 30005 21499 30039
rect 2605 29801 2639 29835
rect 3341 29801 3375 29835
rect 14565 29801 14599 29835
rect 15485 29801 15519 29835
rect 16037 29801 16071 29835
rect 18245 29801 18279 29835
rect 18429 29801 18463 29835
rect 20361 29801 20395 29835
rect 20545 29801 20579 29835
rect 21189 29801 21223 29835
rect 22753 29801 22787 29835
rect 22937 29801 22971 29835
rect 24777 29801 24811 29835
rect 12541 29733 12575 29767
rect 4261 29665 4295 29699
rect 5733 29665 5767 29699
rect 5825 29665 5859 29699
rect 12081 29665 12115 29699
rect 17877 29665 17911 29699
rect 2605 29597 2639 29631
rect 2789 29597 2823 29631
rect 3249 29597 3283 29631
rect 3433 29597 3467 29631
rect 4169 29597 4203 29631
rect 5549 29597 5583 29631
rect 5641 29597 5675 29631
rect 8217 29597 8251 29631
rect 9137 29597 9171 29631
rect 9340 29597 9374 29631
rect 9505 29597 9539 29631
rect 10609 29597 10643 29631
rect 10701 29597 10735 29631
rect 10793 29597 10827 29631
rect 10977 29597 11011 29631
rect 12173 29597 12207 29631
rect 13369 29597 13403 29631
rect 14289 29597 14323 29631
rect 14381 29597 14415 29631
rect 14657 29597 14691 29631
rect 15301 29597 15335 29631
rect 16221 29597 16255 29631
rect 16497 29597 16531 29631
rect 19993 29597 20027 29631
rect 22477 29597 22511 29631
rect 25053 29597 25087 29631
rect 6837 29529 6871 29563
rect 7021 29529 7055 29563
rect 8401 29529 8435 29563
rect 21005 29529 21039 29563
rect 24777 29529 24811 29563
rect 4537 29461 4571 29495
rect 5365 29461 5399 29495
rect 7205 29461 7239 29495
rect 8585 29461 8619 29495
rect 9229 29461 9263 29495
rect 9505 29461 9539 29495
rect 10333 29461 10367 29495
rect 13553 29461 13587 29495
rect 14473 29461 14507 29495
rect 16405 29461 16439 29495
rect 18245 29461 18279 29495
rect 20361 29461 20395 29495
rect 21205 29461 21239 29495
rect 21373 29461 21407 29495
rect 24961 29461 24995 29495
rect 7113 29257 7147 29291
rect 9045 29257 9079 29291
rect 11805 29257 11839 29291
rect 12357 29257 12391 29291
rect 14289 29257 14323 29291
rect 16313 29257 16347 29291
rect 17877 29257 17911 29291
rect 20085 29257 20119 29291
rect 24869 29257 24903 29291
rect 8217 29189 8251 29223
rect 12633 29189 12667 29223
rect 13737 29189 13771 29223
rect 15178 29189 15212 29223
rect 17417 29189 17451 29223
rect 18797 29189 18831 29223
rect 18997 29189 19031 29223
rect 20453 29189 20487 29223
rect 22017 29189 22051 29223
rect 3985 29121 4019 29155
rect 6745 29121 6779 29155
rect 8033 29121 8067 29155
rect 8309 29121 8343 29155
rect 8401 29121 8435 29155
rect 9229 29121 9263 29155
rect 10333 29121 10367 29155
rect 11713 29121 11747 29155
rect 11897 29121 11931 29155
rect 12357 29121 12391 29155
rect 13645 29121 13679 29155
rect 14473 29121 14507 29155
rect 14933 29121 14967 29155
rect 17233 29121 17267 29155
rect 18061 29121 18095 29155
rect 18245 29121 18279 29155
rect 18337 29121 18371 29155
rect 20269 29121 20303 29155
rect 20545 29121 20579 29155
rect 21005 29121 21039 29155
rect 21189 29121 21223 29155
rect 21281 29121 21315 29155
rect 22201 29121 22235 29155
rect 23029 29121 23063 29155
rect 24501 29121 24535 29155
rect 4721 29053 4755 29087
rect 4997 29053 5031 29087
rect 6837 29053 6871 29087
rect 9321 29053 9355 29087
rect 9413 29053 9447 29087
rect 9505 29053 9539 29087
rect 10609 29053 10643 29087
rect 22937 29053 22971 29087
rect 24593 29053 24627 29087
rect 4169 28985 4203 29019
rect 8585 28985 8619 29019
rect 12449 28985 12483 29019
rect 19165 28985 19199 29019
rect 23397 28985 23431 29019
rect 18981 28917 19015 28951
rect 21005 28917 21039 28951
rect 22385 28917 22419 28951
rect 4445 28713 4479 28747
rect 5457 28713 5491 28747
rect 7573 28713 7607 28747
rect 9413 28713 9447 28747
rect 9597 28713 9631 28747
rect 11989 28713 12023 28747
rect 15485 28713 15519 28747
rect 16221 28713 16255 28747
rect 25053 28713 25087 28747
rect 7021 28645 7055 28679
rect 15393 28645 15427 28679
rect 18797 28645 18831 28679
rect 19441 28645 19475 28679
rect 21465 28645 21499 28679
rect 23489 28645 23523 28679
rect 7757 28577 7791 28611
rect 7849 28577 7883 28611
rect 14749 28577 14783 28611
rect 18889 28577 18923 28611
rect 19901 28577 19935 28611
rect 21005 28577 21039 28611
rect 23029 28577 23063 28611
rect 24685 28577 24719 28611
rect 4169 28509 4203 28543
rect 5181 28509 5215 28543
rect 6193 28509 6227 28543
rect 6929 28509 6963 28543
rect 7113 28509 7147 28543
rect 7941 28509 7975 28543
rect 8033 28509 8067 28543
rect 9137 28509 9171 28543
rect 10609 28509 10643 28543
rect 10865 28509 10899 28543
rect 14289 28509 14323 28543
rect 14565 28509 14599 28543
rect 14657 28509 14691 28543
rect 15577 28509 15611 28543
rect 16037 28509 16071 28543
rect 16129 28509 16163 28543
rect 17785 28509 17819 28543
rect 19625 28509 19659 28543
rect 19717 28509 19751 28543
rect 19809 28509 19843 28543
rect 21097 28509 21131 28543
rect 22201 28509 22235 28543
rect 22385 28509 22419 28543
rect 22477 28509 22511 28543
rect 23121 28509 23155 28543
rect 24777 28509 24811 28543
rect 6377 28441 6411 28475
rect 15209 28441 15243 28475
rect 18429 28441 18463 28475
rect 4629 28373 4663 28407
rect 5641 28373 5675 28407
rect 14381 28373 14415 28407
rect 15301 28373 15335 28407
rect 16405 28373 16439 28407
rect 17877 28373 17911 28407
rect 22017 28373 22051 28407
rect 3525 28169 3559 28203
rect 5089 28169 5123 28203
rect 5825 28169 5859 28203
rect 7865 28169 7899 28203
rect 8033 28169 8067 28203
rect 8677 28169 8711 28203
rect 9505 28169 9539 28203
rect 18981 28169 19015 28203
rect 22385 28169 22419 28203
rect 7665 28101 7699 28135
rect 9137 28101 9171 28135
rect 9353 28101 9387 28135
rect 10241 28101 10275 28135
rect 13544 28101 13578 28135
rect 21281 28101 21315 28135
rect 24041 28101 24075 28135
rect 24869 28101 24903 28135
rect 2412 28033 2446 28067
rect 3985 28033 4019 28067
rect 4169 28033 4203 28067
rect 5273 28033 5307 28067
rect 5733 28033 5767 28067
rect 8493 28033 8527 28067
rect 8677 28033 8711 28067
rect 10057 28033 10091 28067
rect 11897 28033 11931 28067
rect 13277 28033 13311 28067
rect 16865 28033 16899 28067
rect 17141 28033 17175 28067
rect 17785 28033 17819 28067
rect 18521 28033 18555 28067
rect 19533 28033 19567 28067
rect 20453 28033 20487 28067
rect 20637 28033 20671 28067
rect 20729 28033 20763 28067
rect 21189 28033 21223 28067
rect 22109 28033 22143 28067
rect 22201 28033 22235 28067
rect 24225 28033 24259 28067
rect 24317 28033 24351 28067
rect 24777 28033 24811 28067
rect 24961 28033 24995 28067
rect 2145 27965 2179 27999
rect 4813 27965 4847 27999
rect 4905 27965 4939 27999
rect 5181 27965 5215 27999
rect 11805 27965 11839 27999
rect 12265 27965 12299 27999
rect 15117 27965 15151 27999
rect 15393 27965 15427 27999
rect 16957 27965 16991 27999
rect 4077 27897 4111 27931
rect 14657 27897 14691 27931
rect 19533 27897 19567 27931
rect 20269 27897 20303 27931
rect 4629 27829 4663 27863
rect 7849 27829 7883 27863
rect 9321 27829 9355 27863
rect 16865 27829 16899 27863
rect 17325 27829 17359 27863
rect 17877 27829 17911 27863
rect 18797 27829 18831 27863
rect 24041 27829 24075 27863
rect 2513 27625 2547 27659
rect 4169 27625 4203 27659
rect 5365 27625 5399 27659
rect 13553 27625 13587 27659
rect 15945 27625 15979 27659
rect 18245 27625 18279 27659
rect 5733 27557 5767 27591
rect 8309 27557 8343 27591
rect 12265 27557 12299 27591
rect 13737 27557 13771 27591
rect 16129 27557 16163 27591
rect 16773 27557 16807 27591
rect 19717 27557 19751 27591
rect 20729 27557 20763 27591
rect 25145 27557 25179 27591
rect 37841 27557 37875 27591
rect 14473 27489 14507 27523
rect 14749 27489 14783 27523
rect 15853 27489 15887 27523
rect 17233 27489 17267 27523
rect 20453 27489 20487 27523
rect 21557 27489 21591 27523
rect 24869 27489 24903 27523
rect 1593 27421 1627 27455
rect 2513 27421 2547 27455
rect 2697 27421 2731 27455
rect 4353 27421 4387 27455
rect 4629 27421 4663 27455
rect 4813 27421 4847 27455
rect 5273 27421 5307 27455
rect 7665 27421 7699 27455
rect 7849 27421 7883 27455
rect 8585 27421 8619 27455
rect 9505 27421 9539 27455
rect 11529 27421 11563 27455
rect 11805 27421 11839 27455
rect 12541 27421 12575 27455
rect 14657 27421 14691 27455
rect 14841 27421 14875 27455
rect 14933 27421 14967 27455
rect 15485 27421 15519 27455
rect 15945 27421 15979 27455
rect 17325 27421 17359 27455
rect 17969 27421 18003 27455
rect 18153 27421 18187 27455
rect 18245 27421 18279 27455
rect 20361 27421 20395 27455
rect 21649 27421 21683 27455
rect 23397 27421 23431 27455
rect 24777 27421 24811 27455
rect 38025 27421 38059 27455
rect 8309 27353 8343 27387
rect 9137 27353 9171 27387
rect 9321 27353 9355 27387
rect 10425 27353 10459 27387
rect 12265 27353 12299 27387
rect 13369 27353 13403 27387
rect 16773 27353 16807 27387
rect 17509 27353 17543 27387
rect 19533 27353 19567 27387
rect 23489 27353 23523 27387
rect 1777 27285 1811 27319
rect 7849 27285 7883 27319
rect 8493 27285 8527 27319
rect 10517 27285 10551 27319
rect 11345 27285 11379 27319
rect 11713 27285 11747 27319
rect 12449 27285 12483 27319
rect 13579 27285 13613 27319
rect 18429 27285 18463 27319
rect 22017 27285 22051 27319
rect 1869 27081 1903 27115
rect 11161 27081 11195 27115
rect 11989 27081 12023 27115
rect 13737 27081 13771 27115
rect 14289 27081 14323 27115
rect 20269 27081 20303 27115
rect 24501 27081 24535 27115
rect 3341 27013 3375 27047
rect 4077 27013 4111 27047
rect 4293 27013 4327 27047
rect 10048 27013 10082 27047
rect 12357 27013 12391 27047
rect 13185 27013 13219 27047
rect 15945 27013 15979 27047
rect 20729 27013 20763 27047
rect 20929 27013 20963 27047
rect 23673 27013 23707 27047
rect 2053 26945 2087 26979
rect 3525 26945 3559 26979
rect 3617 26945 3651 26979
rect 5089 26945 5123 26979
rect 5273 26945 5307 26979
rect 5365 26945 5399 26979
rect 5825 26945 5859 26979
rect 6009 26945 6043 26979
rect 6817 26945 6851 26979
rect 12173 26945 12207 26979
rect 12449 26945 12483 26979
rect 12909 26945 12943 26979
rect 13645 26945 13679 26979
rect 13829 26945 13863 26979
rect 14565 26945 14599 26979
rect 14749 26945 14783 26979
rect 15301 26945 15335 26979
rect 16957 26945 16991 26979
rect 17601 26945 17635 26979
rect 19145 26945 19179 26979
rect 22109 26945 22143 26979
rect 22293 26945 22327 26979
rect 23857 26945 23891 26979
rect 23949 26945 23983 26979
rect 24409 26945 24443 26979
rect 24593 26945 24627 26979
rect 6561 26877 6595 26911
rect 8401 26877 8435 26911
rect 8677 26877 8711 26911
rect 9781 26877 9815 26911
rect 14473 26877 14507 26911
rect 14657 26877 14691 26911
rect 16313 26877 16347 26911
rect 17877 26877 17911 26911
rect 18889 26877 18923 26911
rect 7941 26809 7975 26843
rect 13001 26809 13035 26843
rect 16221 26809 16255 26843
rect 21097 26809 21131 26843
rect 3341 26741 3375 26775
rect 4261 26741 4295 26775
rect 4445 26741 4479 26775
rect 4905 26741 4939 26775
rect 5917 26741 5951 26775
rect 13093 26741 13127 26775
rect 15393 26741 15427 26775
rect 15945 26741 15979 26775
rect 16129 26741 16163 26775
rect 17049 26741 17083 26775
rect 20913 26741 20947 26775
rect 22109 26741 22143 26775
rect 23673 26741 23707 26775
rect 3985 26537 4019 26571
rect 5365 26537 5399 26571
rect 6193 26537 6227 26571
rect 10885 26537 10919 26571
rect 12265 26537 12299 26571
rect 13093 26537 13127 26571
rect 14749 26537 14783 26571
rect 14933 26537 14967 26571
rect 16221 26537 16255 26571
rect 18061 26537 18095 26571
rect 18337 26537 18371 26571
rect 21281 26537 21315 26571
rect 25053 26537 25087 26571
rect 3341 26469 3375 26503
rect 8033 26469 8067 26503
rect 16405 26469 16439 26503
rect 17049 26469 17083 26503
rect 23489 26469 23523 26503
rect 4537 26401 4571 26435
rect 7757 26401 7791 26435
rect 7849 26401 7883 26435
rect 11805 26401 11839 26435
rect 14657 26401 14691 26435
rect 19809 26401 19843 26435
rect 20913 26401 20947 26435
rect 24685 26401 24719 26435
rect 1961 26333 1995 26367
rect 4166 26333 4200 26367
rect 4629 26333 4663 26367
rect 5089 26333 5123 26367
rect 6469 26333 6503 26367
rect 6561 26333 6595 26367
rect 6653 26333 6687 26367
rect 6837 26333 6871 26367
rect 9505 26333 9539 26367
rect 11897 26333 11931 26367
rect 13553 26333 13587 26367
rect 13737 26333 13771 26367
rect 14749 26333 14783 26367
rect 15393 26333 15427 26367
rect 15577 26333 15611 26367
rect 16865 26333 16899 26367
rect 17693 26333 17727 26367
rect 17785 26333 17819 26367
rect 18153 26333 18187 26367
rect 19533 26333 19567 26367
rect 19625 26333 19659 26367
rect 21005 26333 21039 26367
rect 22109 26333 22143 26367
rect 22365 26333 22399 26367
rect 24777 26333 24811 26367
rect 37473 26333 37507 26367
rect 37749 26333 37783 26367
rect 2228 26265 2262 26299
rect 7389 26265 7423 26299
rect 9772 26265 9806 26299
rect 12725 26265 12759 26299
rect 12909 26265 12943 26299
rect 14473 26265 14507 26299
rect 16037 26265 16071 26299
rect 16237 26265 16271 26299
rect 4169 26197 4203 26231
rect 5549 26197 5583 26231
rect 13737 26197 13771 26231
rect 15485 26197 15519 26231
rect 2605 25993 2639 26027
rect 4261 25993 4295 26027
rect 4921 25993 4955 26027
rect 5641 25993 5675 26027
rect 12265 25993 12299 26027
rect 18981 25993 19015 26027
rect 21097 25993 21131 26027
rect 24041 25993 24075 26027
rect 24961 25993 24995 26027
rect 3893 25925 3927 25959
rect 4721 25925 4755 25959
rect 10701 25925 10735 25959
rect 18245 25925 18279 25959
rect 18429 25925 18463 25959
rect 19257 25925 19291 25959
rect 19487 25925 19521 25959
rect 2513 25857 2547 25891
rect 2697 25857 2731 25891
rect 4077 25857 4111 25891
rect 5549 25857 5583 25891
rect 5733 25857 5767 25891
rect 5825 25857 5859 25891
rect 6561 25857 6595 25891
rect 6745 25857 6779 25891
rect 6837 25857 6871 25891
rect 7481 25857 7515 25891
rect 7665 25857 7699 25891
rect 8677 25857 8711 25891
rect 9505 25857 9539 25891
rect 9689 25857 9723 25891
rect 9781 25857 9815 25891
rect 12081 25857 12115 25891
rect 12265 25857 12299 25891
rect 13277 25857 13311 25891
rect 13461 25857 13495 25891
rect 14197 25857 14231 25891
rect 14381 25857 14415 25891
rect 14841 25857 14875 25891
rect 15025 25857 15059 25891
rect 15761 25857 15795 25891
rect 17049 25857 17083 25891
rect 19165 25857 19199 25891
rect 19349 25857 19383 25891
rect 20085 25857 20119 25891
rect 20269 25857 20303 25891
rect 21005 25857 21039 25891
rect 22477 25857 22511 25891
rect 23581 25857 23615 25891
rect 24501 25857 24535 25891
rect 8769 25789 8803 25823
rect 19625 25789 19659 25823
rect 5089 25721 5123 25755
rect 9045 25721 9079 25755
rect 9505 25721 9539 25755
rect 15945 25721 15979 25755
rect 24777 25721 24811 25755
rect 4905 25653 4939 25687
rect 6561 25653 6595 25687
rect 7849 25653 7883 25687
rect 8677 25653 8711 25687
rect 10793 25653 10827 25687
rect 13277 25653 13311 25687
rect 13645 25653 13679 25687
rect 14289 25653 14323 25687
rect 14841 25653 14875 25687
rect 15209 25653 15243 25687
rect 17141 25653 17175 25687
rect 17509 25653 17543 25687
rect 20085 25653 20119 25687
rect 22661 25653 22695 25687
rect 23765 25653 23799 25687
rect 4537 25449 4571 25483
rect 6653 25449 6687 25483
rect 8401 25449 8435 25483
rect 8585 25449 8619 25483
rect 9229 25449 9263 25483
rect 13277 25449 13311 25483
rect 16037 25449 16071 25483
rect 19441 25449 19475 25483
rect 23121 25449 23155 25483
rect 16957 25381 16991 25415
rect 18613 25381 18647 25415
rect 21741 25381 21775 25415
rect 17417 25313 17451 25347
rect 17509 25313 17543 25347
rect 20361 25313 20395 25347
rect 22845 25313 22879 25347
rect 4537 25245 4571 25279
rect 4813 25245 4847 25279
rect 5549 25245 5583 25279
rect 5638 25245 5672 25279
rect 5754 25245 5788 25279
rect 5917 25245 5951 25279
rect 7573 25245 7607 25279
rect 9137 25245 9171 25279
rect 9321 25245 9355 25279
rect 9965 25245 9999 25279
rect 10149 25245 10183 25279
rect 14841 25245 14875 25279
rect 15025 25245 15059 25279
rect 17325 25245 17359 25279
rect 18889 25245 18923 25279
rect 19441 25245 19475 25279
rect 19625 25245 19659 25279
rect 22753 25245 22787 25279
rect 6469 25177 6503 25211
rect 8217 25177 8251 25211
rect 8433 25177 8467 25211
rect 10609 25177 10643 25211
rect 10793 25177 10827 25211
rect 13093 25177 13127 25211
rect 13309 25177 13343 25211
rect 15853 25177 15887 25211
rect 18613 25177 18647 25211
rect 20606 25177 20640 25211
rect 4721 25109 4755 25143
rect 5273 25109 5307 25143
rect 6669 25109 6703 25143
rect 6837 25109 6871 25143
rect 7665 25109 7699 25143
rect 10149 25109 10183 25143
rect 10977 25109 11011 25143
rect 13461 25109 13495 25143
rect 14933 25109 14967 25143
rect 16053 25109 16087 25143
rect 16221 25109 16255 25143
rect 18797 25109 18831 25143
rect 13737 24905 13771 24939
rect 15209 24905 15243 24939
rect 19349 24905 19383 24939
rect 20545 24905 20579 24939
rect 23489 24905 23523 24939
rect 4896 24837 4930 24871
rect 10425 24837 10459 24871
rect 10517 24837 10551 24871
rect 14381 24837 14415 24871
rect 19835 24837 19869 24871
rect 24777 24837 24811 24871
rect 2237 24769 2271 24803
rect 2421 24769 2455 24803
rect 3157 24769 3191 24803
rect 6837 24769 6871 24803
rect 8289 24769 8323 24803
rect 10241 24769 10275 24803
rect 10609 24769 10643 24803
rect 11713 24769 11747 24803
rect 11897 24769 11931 24803
rect 13461 24769 13495 24803
rect 14565 24769 14599 24803
rect 14749 24769 14783 24803
rect 15393 24769 15427 24803
rect 15669 24769 15703 24803
rect 15853 24769 15887 24803
rect 17509 24769 17543 24803
rect 17601 24769 17635 24803
rect 17693 24772 17727 24806
rect 17877 24769 17911 24803
rect 18521 24769 18555 24803
rect 18613 24769 18647 24803
rect 18797 24769 18831 24803
rect 19533 24769 19567 24803
rect 19625 24769 19659 24803
rect 19717 24769 19751 24803
rect 20453 24769 20487 24803
rect 20637 24769 20671 24803
rect 22109 24769 22143 24803
rect 22365 24769 22399 24803
rect 24409 24769 24443 24803
rect 24593 24769 24627 24803
rect 4629 24701 4663 24735
rect 6561 24701 6595 24735
rect 8033 24701 8067 24735
rect 11805 24701 11839 24735
rect 13277 24701 13311 24735
rect 13829 24701 13863 24735
rect 17233 24701 17267 24735
rect 18705 24701 18739 24735
rect 19993 24701 20027 24735
rect 6009 24633 6043 24667
rect 18337 24633 18371 24667
rect 2237 24565 2271 24599
rect 3249 24565 3283 24599
rect 3617 24565 3651 24599
rect 9413 24565 9447 24599
rect 10793 24565 10827 24599
rect 3985 24361 4019 24395
rect 7113 24361 7147 24395
rect 7941 24361 7975 24395
rect 10793 24361 10827 24395
rect 19717 24361 19751 24395
rect 19901 24361 19935 24395
rect 20913 24361 20947 24395
rect 21741 24361 21775 24395
rect 23029 24361 23063 24395
rect 6285 24293 6319 24327
rect 19993 24293 20027 24327
rect 21097 24293 21131 24327
rect 1593 24225 1627 24259
rect 4537 24225 4571 24259
rect 6009 24225 6043 24259
rect 7205 24225 7239 24259
rect 11345 24225 11379 24259
rect 17601 24225 17635 24259
rect 23857 24225 23891 24259
rect 1860 24157 1894 24191
rect 4166 24157 4200 24191
rect 4629 24157 4663 24191
rect 6101 24157 6135 24191
rect 7113 24157 7147 24191
rect 8217 24157 8251 24191
rect 10425 24157 10459 24191
rect 13461 24157 13495 24191
rect 13737 24157 13771 24191
rect 14289 24157 14323 24191
rect 16405 24157 16439 24191
rect 16589 24157 16623 24191
rect 17877 24157 17911 24191
rect 19717 24157 19751 24191
rect 20545 24157 20579 24191
rect 21925 24157 21959 24191
rect 23673 24157 23707 24191
rect 5641 24089 5675 24123
rect 7941 24089 7975 24123
rect 10609 24089 10643 24123
rect 11612 24089 11646 24123
rect 13645 24089 13679 24123
rect 14556 24089 14590 24123
rect 20085 24089 20119 24123
rect 22937 24089 22971 24123
rect 2973 24021 3007 24055
rect 4169 24021 4203 24055
rect 7481 24021 7515 24055
rect 8125 24021 8159 24055
rect 12725 24021 12759 24055
rect 13277 24021 13311 24055
rect 15669 24021 15703 24055
rect 16497 24021 16531 24055
rect 20913 24021 20947 24055
rect 4629 23817 4663 23851
rect 6009 23817 6043 23851
rect 6929 23817 6963 23851
rect 7941 23817 7975 23851
rect 9781 23817 9815 23851
rect 12173 23817 12207 23851
rect 14289 23817 14323 23851
rect 14473 23817 14507 23851
rect 14933 23817 14967 23851
rect 16221 23817 16255 23851
rect 18245 23817 18279 23851
rect 22217 23817 22251 23851
rect 23305 23817 23339 23851
rect 5181 23749 5215 23783
rect 6745 23749 6779 23783
rect 13277 23749 13311 23783
rect 22017 23749 22051 23783
rect 2513 23681 2547 23715
rect 2697 23681 2731 23715
rect 3341 23681 3375 23715
rect 4169 23681 4203 23715
rect 5365 23681 5399 23715
rect 5825 23681 5859 23715
rect 6009 23681 6043 23715
rect 6561 23681 6595 23715
rect 7757 23681 7791 23715
rect 7941 23681 7975 23715
rect 8668 23681 8702 23715
rect 10793 23681 10827 23715
rect 12357 23681 12391 23715
rect 12449 23681 12483 23715
rect 12633 23681 12667 23715
rect 12725 23681 12759 23715
rect 13185 23681 13219 23715
rect 13369 23681 13403 23715
rect 15117 23681 15151 23715
rect 16037 23681 16071 23715
rect 16313 23681 16347 23715
rect 17121 23681 17155 23715
rect 23213 23681 23247 23715
rect 23397 23681 23431 23715
rect 2605 23613 2639 23647
rect 3433 23613 3467 23647
rect 3709 23613 3743 23647
rect 8401 23613 8435 23647
rect 10701 23613 10735 23647
rect 16865 23613 16899 23647
rect 18705 23613 18739 23647
rect 18981 23613 19015 23647
rect 20637 23613 20671 23647
rect 20913 23613 20947 23647
rect 23581 23613 23615 23647
rect 13921 23545 13955 23579
rect 16037 23545 16071 23579
rect 23029 23545 23063 23579
rect 4445 23477 4479 23511
rect 11161 23477 11195 23511
rect 14289 23477 14323 23511
rect 22201 23477 22235 23511
rect 22385 23477 22419 23511
rect 8585 23273 8619 23307
rect 13001 23273 13035 23307
rect 16313 23273 16347 23307
rect 18889 23273 18923 23307
rect 19993 23273 20027 23307
rect 20913 23273 20947 23307
rect 23949 23273 23983 23307
rect 4261 23205 4295 23239
rect 6561 23205 6595 23239
rect 8401 23205 8435 23239
rect 9321 23205 9355 23239
rect 3985 23137 4019 23171
rect 15393 23137 15427 23171
rect 15853 23137 15887 23171
rect 16589 23137 16623 23171
rect 19441 23137 19475 23171
rect 21097 23137 21131 23171
rect 21189 23137 21223 23171
rect 22569 23137 22603 23171
rect 4997 23069 5031 23103
rect 5917 23069 5951 23103
rect 6101 23069 6135 23103
rect 6837 23069 6871 23103
rect 8493 23069 8527 23103
rect 9597 23069 9631 23103
rect 15485 23069 15519 23103
rect 16497 23069 16531 23103
rect 16681 23069 16715 23103
rect 16773 23069 16807 23103
rect 17509 23069 17543 23103
rect 19809 23069 19843 23103
rect 21281 23069 21315 23103
rect 21373 23069 21407 23103
rect 22109 23069 22143 23103
rect 6561 23001 6595 23035
rect 8125 23001 8159 23035
rect 9321 23001 9355 23035
rect 12909 23001 12943 23035
rect 17754 23001 17788 23035
rect 19717 23001 19751 23035
rect 22814 23001 22848 23035
rect 4445 22933 4479 22967
rect 5089 22933 5123 22967
rect 6101 22933 6135 22967
rect 6745 22933 6779 22967
rect 8217 22933 8251 22967
rect 9505 22933 9539 22967
rect 19625 22933 19659 22967
rect 21925 22933 21959 22967
rect 3617 22729 3651 22763
rect 5549 22729 5583 22763
rect 10241 22729 10275 22763
rect 15577 22729 15611 22763
rect 17141 22729 17175 22763
rect 18797 22729 18831 22763
rect 20085 22729 20119 22763
rect 23581 22729 23615 22763
rect 3433 22661 3467 22695
rect 6806 22661 6840 22695
rect 11805 22661 11839 22695
rect 15485 22661 15519 22695
rect 19625 22661 19659 22695
rect 20453 22661 20487 22695
rect 21373 22661 21407 22695
rect 2789 22593 2823 22627
rect 2973 22593 3007 22627
rect 3709 22593 3743 22627
rect 4169 22593 4203 22627
rect 4353 22593 4387 22627
rect 5365 22593 5399 22627
rect 5549 22593 5583 22627
rect 9413 22593 9447 22627
rect 10425 22593 10459 22627
rect 10517 22593 10551 22627
rect 10701 22593 10735 22627
rect 13737 22593 13771 22627
rect 17417 22593 17451 22627
rect 17509 22593 17543 22627
rect 17601 22593 17635 22627
rect 17785 22593 17819 22627
rect 18705 22593 18739 22627
rect 19441 22593 19475 22627
rect 20269 22593 20303 22627
rect 20545 22593 20579 22627
rect 21465 22593 21499 22627
rect 22457 22593 22491 22627
rect 6561 22525 6595 22559
rect 9321 22525 9355 22559
rect 12265 22525 12299 22559
rect 12357 22525 12391 22559
rect 15209 22525 15243 22559
rect 15694 22525 15728 22559
rect 21005 22525 21039 22559
rect 22201 22525 22235 22559
rect 4169 22457 4203 22491
rect 9781 22457 9815 22491
rect 10609 22457 10643 22491
rect 11805 22457 11839 22491
rect 13553 22457 13587 22491
rect 2881 22389 2915 22423
rect 3433 22389 3467 22423
rect 7941 22389 7975 22423
rect 12541 22389 12575 22423
rect 15853 22389 15887 22423
rect 21189 22389 21223 22423
rect 9597 22185 9631 22219
rect 11713 22185 11747 22219
rect 12725 22185 12759 22219
rect 21373 22185 21407 22219
rect 8309 22117 8343 22151
rect 13277 22117 13311 22151
rect 9873 22049 9907 22083
rect 10057 22049 10091 22083
rect 12357 22049 12391 22083
rect 16865 22049 16899 22083
rect 22661 22049 22695 22083
rect 2145 21981 2179 22015
rect 2329 21981 2363 22015
rect 2973 21981 3007 22015
rect 3065 21981 3099 22015
rect 3341 21981 3375 22015
rect 3433 21981 3467 22015
rect 4261 21981 4295 22015
rect 4445 21981 4479 22015
rect 4905 21981 4939 22015
rect 8493 21981 8527 22015
rect 8585 21981 8619 22015
rect 9781 21981 9815 22015
rect 9965 21981 9999 22015
rect 11529 21981 11563 22015
rect 12449 21981 12483 22015
rect 13461 21981 13495 22015
rect 13645 21981 13679 22015
rect 13737 21981 13771 22015
rect 14289 21981 14323 22015
rect 14545 21981 14579 22015
rect 16957 21981 16991 22015
rect 17969 21981 18003 22015
rect 18061 21981 18095 22015
rect 18705 21981 18739 22015
rect 18889 21981 18923 22015
rect 19441 21981 19475 22015
rect 21557 21981 21591 22015
rect 21741 21981 21775 22015
rect 21833 21981 21867 22015
rect 22385 21981 22419 22015
rect 2237 21913 2271 21947
rect 3157 21913 3191 21947
rect 4353 21913 4387 21947
rect 5150 21913 5184 21947
rect 8309 21913 8343 21947
rect 11161 21913 11195 21947
rect 11437 21913 11471 21947
rect 17785 21913 17819 21947
rect 18797 21913 18831 21947
rect 19686 21913 19720 21947
rect 2789 21845 2823 21879
rect 6285 21845 6319 21879
rect 11345 21845 11379 21879
rect 15669 21845 15703 21879
rect 17325 21845 17359 21879
rect 17883 21845 17917 21879
rect 20821 21845 20855 21879
rect 2789 21641 2823 21675
rect 4353 21641 4387 21675
rect 7389 21641 7423 21675
rect 9781 21641 9815 21675
rect 14933 21641 14967 21675
rect 19809 21641 19843 21675
rect 21097 21641 21131 21675
rect 23857 21641 23891 21675
rect 2421 21573 2455 21607
rect 6745 21573 6779 21607
rect 20821 21573 20855 21607
rect 21005 21573 21039 21607
rect 2605 21505 2639 21539
rect 3433 21505 3467 21539
rect 4537 21505 4571 21539
rect 4629 21505 4663 21539
rect 4905 21505 4939 21539
rect 5641 21505 5675 21539
rect 6653 21505 6687 21539
rect 7573 21505 7607 21539
rect 7849 21505 7883 21539
rect 8401 21505 8435 21539
rect 8585 21505 8619 21539
rect 8677 21505 8711 21539
rect 8861 21505 8895 21539
rect 8953 21505 8987 21539
rect 9597 21505 9631 21539
rect 10701 21505 10735 21539
rect 10977 21505 11011 21539
rect 12265 21505 12299 21539
rect 15209 21505 15243 21539
rect 15669 21505 15703 21539
rect 17141 21505 17175 21539
rect 17408 21505 17442 21539
rect 19533 21505 19567 21539
rect 19625 21505 19659 21539
rect 21097 21505 21131 21539
rect 22744 21505 22778 21539
rect 3341 21437 3375 21471
rect 4813 21437 4847 21471
rect 5733 21437 5767 21471
rect 7665 21437 7699 21471
rect 9413 21437 9447 21471
rect 10793 21437 10827 21471
rect 12173 21437 12207 21471
rect 15485 21437 15519 21471
rect 22477 21437 22511 21471
rect 3801 21369 3835 21403
rect 6009 21369 6043 21403
rect 7757 21369 7791 21403
rect 12633 21369 12667 21403
rect 10977 21301 11011 21335
rect 11161 21301 11195 21335
rect 15301 21301 15335 21335
rect 15393 21301 15427 21335
rect 18521 21301 18555 21335
rect 6837 21097 6871 21131
rect 7113 21097 7147 21131
rect 7941 21097 7975 21131
rect 9597 21097 9631 21131
rect 10425 21097 10459 21131
rect 10793 21097 10827 21131
rect 13461 21097 13495 21131
rect 15393 21097 15427 21131
rect 16681 21097 16715 21131
rect 17693 21097 17727 21131
rect 19717 21097 19751 21131
rect 21465 21097 21499 21131
rect 23029 21097 23063 21131
rect 2329 21029 2363 21063
rect 5825 21029 5859 21063
rect 10701 21029 10735 21063
rect 12357 21029 12391 21063
rect 19625 21029 19659 21063
rect 22385 21029 22419 21063
rect 5549 20961 5583 20995
rect 6837 20961 6871 20995
rect 9229 20961 9263 20995
rect 10885 20961 10919 20995
rect 11897 20961 11931 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 19809 20961 19843 20995
rect 22109 20961 22143 20995
rect 22569 20961 22603 20995
rect 1593 20893 1627 20927
rect 2513 20893 2547 20927
rect 3249 20893 3283 20927
rect 3433 20893 3467 20927
rect 5733 20893 5767 20927
rect 5917 20893 5951 20927
rect 6009 20893 6043 20927
rect 6561 20893 6595 20927
rect 8125 20893 8159 20927
rect 8309 20893 8343 20927
rect 8401 20893 8435 20927
rect 9321 20893 9355 20927
rect 10977 20893 11011 20927
rect 11161 20893 11195 20927
rect 11621 20893 11655 20927
rect 11713 20893 11747 20927
rect 12357 20893 12391 20927
rect 12541 20893 12575 20927
rect 15577 20893 15611 20927
rect 15853 20893 15887 20927
rect 17969 20893 18003 20927
rect 18521 20893 18555 20927
rect 19533 20893 19567 20927
rect 21097 20893 21131 20927
rect 23213 20893 23247 20927
rect 4445 20825 4479 20859
rect 4629 20825 4663 20859
rect 13369 20825 13403 20859
rect 15761 20825 15795 20859
rect 16313 20825 16347 20859
rect 16497 20825 16531 20859
rect 17693 20825 17727 20859
rect 18797 20825 18831 20859
rect 1777 20757 1811 20791
rect 3433 20757 3467 20791
rect 11897 20757 11931 20791
rect 17877 20757 17911 20791
rect 21465 20757 21499 20791
rect 21649 20757 21683 20791
rect 6929 20553 6963 20587
rect 9705 20553 9739 20587
rect 10701 20553 10735 20587
rect 11713 20553 11747 20587
rect 14289 20553 14323 20587
rect 20193 20553 20227 20587
rect 20821 20553 20855 20587
rect 9505 20485 9539 20519
rect 19993 20485 20027 20519
rect 2145 20417 2179 20451
rect 2329 20417 2363 20451
rect 3157 20417 3191 20451
rect 4077 20417 4111 20451
rect 4261 20417 4295 20451
rect 5549 20417 5583 20451
rect 5825 20417 5859 20451
rect 6009 20417 6043 20451
rect 7113 20417 7147 20451
rect 7389 20417 7423 20451
rect 7573 20417 7607 20451
rect 10885 20417 10919 20451
rect 11161 20417 11195 20451
rect 11897 20417 11931 20451
rect 12173 20417 12207 20451
rect 12909 20417 12943 20451
rect 14565 20417 14599 20451
rect 14749 20417 14783 20451
rect 15577 20417 15611 20451
rect 15761 20417 15795 20451
rect 15945 20417 15979 20451
rect 16313 20417 16347 20451
rect 17785 20417 17819 20451
rect 18521 20417 18555 20451
rect 18705 20417 18739 20451
rect 19165 20417 19199 20451
rect 19257 20417 19291 20451
rect 21005 20417 21039 20451
rect 21281 20417 21315 20451
rect 22109 20417 22143 20451
rect 22937 20417 22971 20451
rect 3433 20349 3467 20383
rect 4353 20349 4387 20383
rect 12081 20349 12115 20383
rect 13001 20349 13035 20383
rect 14473 20349 14507 20383
rect 14657 20349 14691 20383
rect 21097 20349 21131 20383
rect 21189 20349 21223 20383
rect 3341 20281 3375 20315
rect 9873 20281 9907 20315
rect 11989 20281 12023 20315
rect 17969 20281 18003 20315
rect 2145 20213 2179 20247
rect 3249 20213 3283 20247
rect 3893 20213 3927 20247
rect 5365 20213 5399 20247
rect 9689 20213 9723 20247
rect 11069 20213 11103 20247
rect 13277 20213 13311 20247
rect 15577 20213 15611 20247
rect 18613 20213 18647 20247
rect 19349 20213 19383 20247
rect 19533 20213 19567 20247
rect 20177 20213 20211 20247
rect 20361 20213 20395 20247
rect 22201 20213 22235 20247
rect 22753 20213 22787 20247
rect 3985 20009 4019 20043
rect 4537 20009 4571 20043
rect 5641 20009 5675 20043
rect 6377 20009 6411 20043
rect 6837 20009 6871 20043
rect 8309 20009 8343 20043
rect 11989 20009 12023 20043
rect 16129 20009 16163 20043
rect 18337 20009 18371 20043
rect 19901 20009 19935 20043
rect 21281 20009 21315 20043
rect 23397 20009 23431 20043
rect 2973 19941 3007 19975
rect 8493 19941 8527 19975
rect 11529 19941 11563 19975
rect 14933 19941 14967 19975
rect 16221 19941 16255 19975
rect 20085 19941 20119 19975
rect 6469 19873 6503 19907
rect 9413 19873 9447 19907
rect 11069 19873 11103 19907
rect 15393 19873 15427 19907
rect 16405 19873 16439 19907
rect 16957 19873 16991 19907
rect 19717 19873 19751 19907
rect 20913 19873 20947 19907
rect 1593 19805 1627 19839
rect 1860 19805 1894 19839
rect 4110 19805 4144 19839
rect 4629 19805 4663 19839
rect 6377 19805 6411 19839
rect 6653 19805 6687 19839
rect 7297 19805 7331 19839
rect 7481 19805 7515 19839
rect 9137 19805 9171 19839
rect 11161 19805 11195 19839
rect 11989 19805 12023 19839
rect 12173 19805 12207 19839
rect 13093 19805 13127 19839
rect 13241 19805 13275 19839
rect 13599 19805 13633 19839
rect 15485 19805 15519 19839
rect 15669 19805 15703 19839
rect 16129 19805 16163 19839
rect 19441 19805 19475 19839
rect 19901 19805 19935 19839
rect 21097 19805 21131 19839
rect 22017 19805 22051 19839
rect 22284 19805 22318 19839
rect 5549 19737 5583 19771
rect 7389 19737 7423 19771
rect 8125 19737 8159 19771
rect 8325 19737 8359 19771
rect 13369 19737 13403 19771
rect 13461 19737 13495 19771
rect 14933 19737 14967 19771
rect 17224 19737 17258 19771
rect 4169 19669 4203 19703
rect 13737 19669 13771 19703
rect 3525 19465 3559 19499
rect 5365 19465 5399 19499
rect 14841 19465 14875 19499
rect 16037 19465 16071 19499
rect 16313 19465 16347 19499
rect 18061 19465 18095 19499
rect 20729 19465 20763 19499
rect 1685 19397 1719 19431
rect 4353 19397 4387 19431
rect 4569 19397 4603 19431
rect 18981 19397 19015 19431
rect 20361 19397 20395 19431
rect 20577 19397 20611 19431
rect 21465 19397 21499 19431
rect 3157 19329 3191 19363
rect 5273 19329 5307 19363
rect 6561 19329 6595 19363
rect 6745 19329 6779 19363
rect 7481 19329 7515 19363
rect 8585 19329 8619 19363
rect 8769 19329 8803 19363
rect 9505 19329 9539 19363
rect 10885 19329 10919 19363
rect 11069 19329 11103 19363
rect 12817 19329 12851 19363
rect 13277 19329 13311 19363
rect 13461 19329 13495 19363
rect 13553 19329 13587 19363
rect 13829 19329 13863 19363
rect 15025 19329 15059 19363
rect 15945 19329 15979 19363
rect 16129 19329 16163 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 18153 19329 18187 19363
rect 18705 19329 18739 19363
rect 19441 19329 19475 19363
rect 19625 19329 19659 19363
rect 21189 19329 21223 19363
rect 22017 19329 22051 19363
rect 22201 19329 22235 19363
rect 3065 19261 3099 19295
rect 8861 19261 8895 19295
rect 9413 19261 9447 19295
rect 13737 19261 13771 19295
rect 15301 19261 15335 19295
rect 15761 19261 15795 19295
rect 17693 19261 17727 19295
rect 18981 19261 19015 19295
rect 21281 19261 21315 19295
rect 21465 19261 21499 19295
rect 1869 19193 1903 19227
rect 4721 19193 4755 19227
rect 10885 19193 10919 19227
rect 15209 19193 15243 19227
rect 16865 19193 16899 19227
rect 18797 19193 18831 19227
rect 4537 19125 4571 19159
rect 6561 19125 6595 19159
rect 6929 19125 6963 19159
rect 7573 19125 7607 19159
rect 7941 19125 7975 19159
rect 8401 19125 8435 19159
rect 9781 19125 9815 19159
rect 12633 19125 12667 19159
rect 13645 19125 13679 19159
rect 17877 19125 17911 19159
rect 19809 19125 19843 19159
rect 20545 19125 20579 19159
rect 22017 19125 22051 19159
rect 38301 19125 38335 19159
rect 3341 18921 3375 18955
rect 5641 18921 5675 18955
rect 6469 18921 6503 18955
rect 8401 18921 8435 18955
rect 8585 18921 8619 18955
rect 14289 18921 14323 18955
rect 14749 18921 14783 18955
rect 17693 18921 17727 18955
rect 18705 18921 18739 18955
rect 19625 18921 19659 18955
rect 22569 18921 22603 18955
rect 9367 18853 9401 18887
rect 11069 18853 11103 18887
rect 12725 18853 12759 18887
rect 16037 18853 16071 18887
rect 5825 18785 5859 18819
rect 7481 18785 7515 18819
rect 10609 18785 10643 18819
rect 18061 18785 18095 18819
rect 3249 18717 3283 18751
rect 4445 18717 4479 18751
rect 4537 18717 4571 18751
rect 5549 18717 5583 18751
rect 7573 18717 7607 18751
rect 9137 18717 9171 18751
rect 10701 18717 10735 18751
rect 12541 18717 12575 18751
rect 14473 18717 14507 18751
rect 14565 18717 14599 18751
rect 15853 18717 15887 18751
rect 17877 18717 17911 18751
rect 18153 18717 18187 18751
rect 18613 18717 18647 18751
rect 20177 18717 20211 18751
rect 20361 18717 20395 18751
rect 21189 18717 21223 18751
rect 21456 18717 21490 18751
rect 6285 18649 6319 18683
rect 8217 18649 8251 18683
rect 13369 18649 13403 18683
rect 14289 18649 14323 18683
rect 17049 18649 17083 18683
rect 19533 18649 19567 18683
rect 4721 18581 4755 18615
rect 5825 18581 5859 18615
rect 6485 18581 6519 18615
rect 6653 18581 6687 18615
rect 7113 18581 7147 18615
rect 7757 18581 7791 18615
rect 8427 18581 8461 18615
rect 13461 18581 13495 18615
rect 17141 18581 17175 18615
rect 20269 18581 20303 18615
rect 3893 18377 3927 18411
rect 6929 18377 6963 18411
rect 10149 18377 10183 18411
rect 10793 18377 10827 18411
rect 14105 18377 14139 18411
rect 18429 18377 18463 18411
rect 20729 18377 20763 18411
rect 3249 18309 3283 18343
rect 5733 18309 5767 18343
rect 6561 18309 6595 18343
rect 6777 18309 6811 18343
rect 9014 18309 9048 18343
rect 10701 18309 10735 18343
rect 12817 18309 12851 18343
rect 17785 18309 17819 18343
rect 19616 18309 19650 18343
rect 2973 18241 3007 18275
rect 3893 18241 3927 18275
rect 4629 18241 4663 18275
rect 4721 18241 4755 18275
rect 4997 18241 5031 18275
rect 5549 18241 5583 18275
rect 7849 18241 7883 18275
rect 8033 18241 8067 18275
rect 8125 18241 8159 18275
rect 11897 18241 11931 18275
rect 12081 18241 12115 18275
rect 12633 18241 12667 18275
rect 13461 18241 13495 18275
rect 13554 18241 13588 18275
rect 13737 18241 13771 18275
rect 13829 18241 13863 18275
rect 13967 18241 14001 18275
rect 15209 18241 15243 18275
rect 17601 18241 17635 18275
rect 18337 18241 18371 18275
rect 19349 18241 19383 18275
rect 3065 18173 3099 18207
rect 3249 18173 3283 18207
rect 4905 18173 4939 18207
rect 7941 18173 7975 18207
rect 8769 18173 8803 18207
rect 12173 18173 12207 18207
rect 15301 18173 15335 18207
rect 15577 18173 15611 18207
rect 4445 18037 4479 18071
rect 6745 18037 6779 18071
rect 7665 18037 7699 18071
rect 11713 18037 11747 18071
rect 13001 18037 13035 18071
rect 4537 17833 4571 17867
rect 7757 17833 7791 17867
rect 12449 17833 12483 17867
rect 12633 17833 12667 17867
rect 13093 17833 13127 17867
rect 15301 17833 15335 17867
rect 17969 17833 18003 17867
rect 18613 17833 18647 17867
rect 6469 17765 6503 17799
rect 13553 17765 13587 17799
rect 15853 17765 15887 17799
rect 4261 17697 4295 17731
rect 6193 17697 6227 17731
rect 10057 17697 10091 17731
rect 11529 17697 11563 17731
rect 15117 17697 15151 17731
rect 16221 17697 16255 17731
rect 17693 17697 17727 17731
rect 3249 17629 3283 17663
rect 4169 17629 4203 17663
rect 4997 17629 5031 17663
rect 5181 17629 5215 17663
rect 6101 17629 6135 17663
rect 7353 17629 7387 17663
rect 7471 17623 7505 17657
rect 7573 17623 7607 17657
rect 10241 17629 10275 17663
rect 11253 17629 11287 17663
rect 13277 17629 13311 17663
rect 13369 17629 13403 17663
rect 13645 17629 13679 17663
rect 15025 17629 15059 17663
rect 16037 17629 16071 17663
rect 16129 17629 16163 17663
rect 16313 17629 16347 17663
rect 17601 17629 17635 17663
rect 3433 17561 3467 17595
rect 11345 17561 11379 17595
rect 12265 17561 12299 17595
rect 18429 17561 18463 17595
rect 5365 17493 5399 17527
rect 10425 17493 10459 17527
rect 10885 17493 10919 17527
rect 12465 17493 12499 17527
rect 18629 17493 18663 17527
rect 18797 17493 18831 17527
rect 4813 17289 4847 17323
rect 7113 17289 7147 17323
rect 19901 17289 19935 17323
rect 5365 17221 5399 17255
rect 10793 17221 10827 17255
rect 3700 17153 3734 17187
rect 6745 17153 6779 17187
rect 7849 17153 7883 17187
rect 9321 17153 9355 17187
rect 9505 17153 9539 17187
rect 10149 17153 10183 17187
rect 10977 17153 11011 17187
rect 12449 17153 12483 17187
rect 12705 17153 12739 17187
rect 14473 17153 14507 17187
rect 14657 17153 14691 17187
rect 15117 17153 15151 17187
rect 15301 17153 15335 17187
rect 15393 17153 15427 17187
rect 15521 17153 15555 17187
rect 16037 17153 16071 17187
rect 16221 17153 16255 17187
rect 17509 17153 17543 17187
rect 18777 17153 18811 17187
rect 3433 17085 3467 17119
rect 6837 17085 6871 17119
rect 7665 17085 7699 17119
rect 9137 17085 9171 17119
rect 11161 17085 11195 17119
rect 15209 17085 15243 17119
rect 18521 17085 18555 17119
rect 5549 17017 5583 17051
rect 17693 17017 17727 17051
rect 8033 16949 8067 16983
rect 9965 16949 9999 16983
rect 13829 16949 13863 16983
rect 14473 16949 14507 16983
rect 16129 16949 16163 16983
rect 4077 16745 4111 16779
rect 8401 16745 8435 16779
rect 11161 16745 11195 16779
rect 15025 16745 15059 16779
rect 15945 16745 15979 16779
rect 18337 16745 18371 16779
rect 12909 16677 12943 16711
rect 16497 16677 16531 16711
rect 7021 16609 7055 16643
rect 9137 16609 9171 16643
rect 11805 16609 11839 16643
rect 12449 16609 12483 16643
rect 14933 16609 14967 16643
rect 15577 16609 15611 16643
rect 17601 16609 17635 16643
rect 17693 16609 17727 16643
rect 17877 16609 17911 16643
rect 4261 16541 4295 16575
rect 6561 16541 6595 16575
rect 9404 16541 9438 16575
rect 12541 16541 12575 16575
rect 13369 16541 13403 16575
rect 13461 16541 13495 16575
rect 14841 16541 14875 16575
rect 15761 16541 15795 16575
rect 16405 16541 16439 16575
rect 16589 16541 16623 16575
rect 18521 16541 18555 16575
rect 7288 16473 7322 16507
rect 11529 16473 11563 16507
rect 15117 16473 15151 16507
rect 6377 16405 6411 16439
rect 10517 16405 10551 16439
rect 11621 16405 11655 16439
rect 17233 16405 17267 16439
rect 7205 16201 7239 16235
rect 10333 16201 10367 16235
rect 11069 16201 11103 16235
rect 14933 16201 14967 16235
rect 17233 16201 17267 16235
rect 19073 16201 19107 16235
rect 10977 16133 11011 16167
rect 15945 16133 15979 16167
rect 16865 16133 16899 16167
rect 17065 16133 17099 16167
rect 7389 16065 7423 16099
rect 9045 16065 9079 16099
rect 10149 16065 10183 16099
rect 10425 16065 10459 16099
rect 11897 16065 11931 16099
rect 11989 16065 12023 16099
rect 12265 16065 12299 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 13737 16065 13771 16099
rect 15117 16065 15151 16099
rect 15301 16065 15335 16099
rect 15853 16065 15887 16099
rect 18981 16065 19015 16099
rect 13553 15997 13587 16031
rect 15393 15997 15427 16031
rect 16221 15997 16255 16031
rect 17693 15997 17727 16031
rect 17969 15997 18003 16031
rect 10149 15929 10183 15963
rect 9229 15861 9263 15895
rect 11713 15861 11747 15895
rect 12173 15861 12207 15895
rect 12817 15861 12851 15895
rect 13093 15861 13127 15895
rect 13921 15861 13955 15895
rect 16129 15861 16163 15895
rect 16313 15861 16347 15895
rect 17049 15861 17083 15895
rect 11345 15657 11379 15691
rect 14841 15657 14875 15691
rect 18797 15657 18831 15691
rect 12633 15589 12667 15623
rect 15393 15589 15427 15623
rect 9321 15521 9355 15555
rect 11529 15521 11563 15555
rect 11704 15521 11738 15555
rect 11805 15521 11839 15555
rect 15485 15521 15519 15555
rect 16865 15521 16899 15555
rect 9137 15453 9171 15487
rect 10057 15453 10091 15487
rect 10333 15453 10367 15487
rect 11610 15453 11644 15487
rect 12909 15453 12943 15487
rect 13001 15453 13035 15487
rect 15022 15453 15056 15487
rect 16497 15453 16531 15487
rect 16589 15453 16623 15487
rect 16957 15453 16991 15487
rect 17417 15453 17451 15487
rect 19441 15453 19475 15487
rect 19625 15453 19659 15487
rect 12817 15385 12851 15419
rect 16221 15385 16255 15419
rect 17684 15385 17718 15419
rect 19533 15385 19567 15419
rect 13185 15317 13219 15351
rect 15025 15317 15059 15351
rect 16681 15317 16715 15351
rect 9781 15113 9815 15147
rect 10425 15113 10459 15147
rect 11713 15113 11747 15147
rect 13369 15113 13403 15147
rect 15025 15113 15059 15147
rect 17233 15113 17267 15147
rect 17049 15045 17083 15079
rect 8401 14977 8435 15011
rect 8668 14977 8702 15011
rect 10366 14977 10400 15011
rect 10885 14977 10919 15011
rect 12081 14977 12115 15011
rect 12173 14977 12207 15011
rect 13001 14977 13035 15011
rect 13093 14977 13127 15011
rect 14197 14977 14231 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 14565 14977 14599 15011
rect 15301 14977 15335 15011
rect 16865 14977 16899 15011
rect 17693 14977 17727 15011
rect 15209 14909 15243 14943
rect 15393 14909 15427 14943
rect 15485 14909 15519 14943
rect 17969 14909 18003 14943
rect 10793 14841 10827 14875
rect 10241 14773 10275 14807
rect 12357 14773 12391 14807
rect 13185 14773 13219 14807
rect 14013 14773 14047 14807
rect 9137 14569 9171 14603
rect 10885 14569 10919 14603
rect 11897 14569 11931 14603
rect 12541 14569 12575 14603
rect 12633 14569 12667 14603
rect 13645 14569 13679 14603
rect 14473 14569 14507 14603
rect 17049 14569 17083 14603
rect 17141 14569 17175 14603
rect 17969 14569 18003 14603
rect 17877 14501 17911 14535
rect 11069 14433 11103 14467
rect 12725 14433 12759 14467
rect 18061 14433 18095 14467
rect 18153 14433 18187 14467
rect 9137 14365 9171 14399
rect 9321 14365 9355 14399
rect 10793 14365 10827 14399
rect 11529 14365 11563 14399
rect 11713 14365 11747 14399
rect 12449 14365 12483 14399
rect 13369 14365 13403 14399
rect 13461 14365 13495 14399
rect 13737 14365 13771 14399
rect 14381 14365 14415 14399
rect 15025 14365 15059 14399
rect 15301 14365 15335 14399
rect 16865 14365 16899 14399
rect 16957 14365 16991 14399
rect 17325 14365 17359 14399
rect 17785 14365 17819 14399
rect 19625 14365 19659 14399
rect 11069 14297 11103 14331
rect 13185 14229 13219 14263
rect 16589 14229 16623 14263
rect 19441 14229 19475 14263
rect 12265 14025 12299 14059
rect 15117 14025 15151 14059
rect 15485 14025 15519 14059
rect 18521 14025 18555 14059
rect 9597 13957 9631 13991
rect 16313 13957 16347 13991
rect 1593 13889 1627 13923
rect 9781 13889 9815 13923
rect 9873 13889 9907 13923
rect 10517 13889 10551 13923
rect 12262 13889 12296 13923
rect 12725 13889 12759 13923
rect 13553 13889 13587 13923
rect 13829 13889 13863 13923
rect 15301 13889 15335 13923
rect 15577 13889 15611 13923
rect 16129 13889 16163 13923
rect 17141 13889 17175 13923
rect 17397 13889 17431 13923
rect 10609 13821 10643 13855
rect 12633 13753 12667 13787
rect 1777 13685 1811 13719
rect 9597 13685 9631 13719
rect 10885 13685 10919 13719
rect 12081 13685 12115 13719
rect 10885 13481 10919 13515
rect 13645 13481 13679 13515
rect 15117 13481 15151 13515
rect 17049 13481 17083 13515
rect 9505 13345 9539 13379
rect 11621 13277 11655 13311
rect 11805 13277 11839 13311
rect 12265 13277 12299 13311
rect 14933 13277 14967 13311
rect 15669 13277 15703 13311
rect 15936 13277 15970 13311
rect 9772 13209 9806 13243
rect 11713 13209 11747 13243
rect 12510 13209 12544 13243
rect 14749 13209 14783 13243
rect 9965 12937 9999 12971
rect 10885 12937 10919 12971
rect 13277 12937 13311 12971
rect 14197 12937 14231 12971
rect 15485 12937 15519 12971
rect 18613 12937 18647 12971
rect 15301 12869 15335 12903
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 13185 12801 13219 12835
rect 13369 12801 13403 12835
rect 13829 12801 13863 12835
rect 14013 12801 14047 12835
rect 14657 12801 14691 12835
rect 14841 12801 14875 12835
rect 15577 12801 15611 12835
rect 18521 12801 18555 12835
rect 38301 12801 38335 12835
rect 14749 12665 14783 12699
rect 15301 12665 15335 12699
rect 38117 12597 38151 12631
rect 17509 12393 17543 12427
rect 17325 12325 17359 12359
rect 17049 12257 17083 12291
rect 1593 7361 1627 7395
rect 1777 7157 1811 7191
rect 1777 6953 1811 6987
rect 1961 6749 1995 6783
rect 37381 5797 37415 5831
rect 37565 5661 37599 5695
rect 38025 5661 38059 5695
rect 38209 5525 38243 5559
rect 25605 3009 25639 3043
rect 32505 3009 32539 3043
rect 32781 3009 32815 3043
rect 25237 2873 25271 2907
rect 25789 2805 25823 2839
rect 32321 2805 32355 2839
rect 6561 2601 6595 2635
rect 19441 2601 19475 2635
rect 1869 2465 1903 2499
rect 1593 2397 1627 2431
rect 6745 2397 6779 2431
rect 13001 2397 13035 2431
rect 19625 2397 19659 2431
rect 25881 2397 25915 2431
rect 32321 2397 32355 2431
rect 38025 2397 38059 2431
rect 13185 2261 13219 2295
rect 26065 2261 26099 2295
rect 32505 2261 32539 2295
rect 38209 2261 38243 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 7098 37272 7104 37324
rect 7156 37312 7162 37324
rect 7193 37315 7251 37321
rect 7193 37312 7205 37315
rect 7156 37284 7205 37312
rect 7156 37272 7162 37284
rect 7193 37281 7205 37284
rect 7239 37281 7251 37315
rect 7193 37275 7251 37281
rect 658 37204 664 37256
rect 716 37244 722 37256
rect 1765 37247 1823 37253
rect 1765 37244 1777 37247
rect 716 37216 1777 37244
rect 716 37204 722 37216
rect 1765 37213 1777 37216
rect 1811 37213 1823 37247
rect 7469 37247 7527 37253
rect 7469 37244 7481 37247
rect 1765 37207 1823 37213
rect 7116 37216 7481 37244
rect 7116 37188 7144 37216
rect 7469 37213 7481 37216
rect 7515 37213 7527 37247
rect 7469 37207 7527 37213
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37244 14335 37247
rect 19426 37244 19432 37256
rect 14323 37216 19432 37244
rect 14323 37213 14335 37216
rect 14277 37207 14335 37213
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 19978 37204 19984 37256
rect 20036 37244 20042 37256
rect 20257 37247 20315 37253
rect 20257 37244 20269 37247
rect 20036 37216 20269 37244
rect 20036 37204 20042 37216
rect 20257 37213 20269 37216
rect 20303 37213 20315 37247
rect 27154 37244 27160 37256
rect 27115 37216 27160 37244
rect 20257 37207 20315 37213
rect 27154 37204 27160 37216
rect 27212 37204 27218 37256
rect 32950 37244 32956 37256
rect 32911 37216 32956 37244
rect 32950 37204 32956 37216
rect 33008 37204 33014 37256
rect 37826 37204 37832 37256
rect 37884 37244 37890 37256
rect 38013 37247 38071 37253
rect 38013 37244 38025 37247
rect 37884 37216 38025 37244
rect 37884 37204 37890 37216
rect 38013 37213 38025 37216
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 7098 37136 7104 37188
rect 7156 37136 7162 37188
rect 1581 37111 1639 37117
rect 1581 37077 1593 37111
rect 1627 37108 1639 37111
rect 3786 37108 3792 37120
rect 1627 37080 3792 37108
rect 1627 37077 1639 37080
rect 1581 37071 1639 37077
rect 3786 37068 3792 37080
rect 3844 37068 3850 37120
rect 13814 37068 13820 37120
rect 13872 37108 13878 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 13872 37080 14473 37108
rect 13872 37068 13878 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 20070 37108 20076 37120
rect 20031 37080 20076 37108
rect 14461 37071 14519 37077
rect 20070 37068 20076 37080
rect 20128 37068 20134 37120
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 26476 37080 27353 37108
rect 26476 37068 26482 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 32858 37068 32864 37120
rect 32916 37108 32922 37120
rect 33137 37111 33195 37117
rect 33137 37108 33149 37111
rect 32916 37080 33149 37108
rect 32916 37068 32922 37080
rect 33137 37077 33149 37080
rect 33183 37077 33195 37111
rect 33137 37071 33195 37077
rect 38197 37111 38255 37117
rect 38197 37077 38209 37111
rect 38243 37108 38255 37111
rect 39298 37108 39304 37120
rect 38243 37080 39304 37108
rect 38243 37077 38255 37080
rect 38197 37071 38255 37077
rect 39298 37068 39304 37080
rect 39356 37068 39362 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 19426 36904 19432 36916
rect 19387 36876 19432 36904
rect 19426 36864 19432 36876
rect 19484 36864 19490 36916
rect 19613 36771 19671 36777
rect 19613 36737 19625 36771
rect 19659 36768 19671 36771
rect 20070 36768 20076 36780
rect 19659 36740 20076 36768
rect 19659 36737 19671 36740
rect 19613 36731 19671 36737
rect 20070 36728 20076 36740
rect 20128 36728 20134 36780
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1581 34595 1639 34601
rect 1581 34561 1593 34595
rect 1627 34592 1639 34595
rect 1670 34592 1676 34604
rect 1627 34564 1676 34592
rect 1627 34561 1639 34564
rect 1581 34555 1639 34561
rect 1670 34552 1676 34564
rect 1728 34552 1734 34604
rect 1762 34388 1768 34400
rect 1723 34360 1768 34388
rect 1762 34348 1768 34360
rect 1820 34348 1826 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 17310 34116 17316 34128
rect 13740 34088 17316 34116
rect 9858 33980 9864 33992
rect 9819 33952 9864 33980
rect 9858 33940 9864 33952
rect 9916 33940 9922 33992
rect 12345 33983 12403 33989
rect 12345 33949 12357 33983
rect 12391 33980 12403 33983
rect 12618 33980 12624 33992
rect 12391 33952 12624 33980
rect 12391 33949 12403 33952
rect 12345 33943 12403 33949
rect 12618 33940 12624 33952
rect 12676 33980 12682 33992
rect 13740 33989 13768 34088
rect 17310 34076 17316 34088
rect 17368 34076 17374 34128
rect 13906 34008 13912 34060
rect 13964 34048 13970 34060
rect 14645 34051 14703 34057
rect 14645 34048 14657 34051
rect 13964 34020 14657 34048
rect 13964 34008 13970 34020
rect 14645 34017 14657 34020
rect 14691 34048 14703 34051
rect 16206 34048 16212 34060
rect 14691 34020 16212 34048
rect 14691 34017 14703 34020
rect 14645 34011 14703 34017
rect 16206 34008 16212 34020
rect 16264 34008 16270 34060
rect 13725 33983 13783 33989
rect 13725 33980 13737 33983
rect 12676 33952 13737 33980
rect 12676 33940 12682 33952
rect 13725 33949 13737 33952
rect 13771 33949 13783 33983
rect 14366 33980 14372 33992
rect 14327 33952 14372 33980
rect 13725 33943 13783 33949
rect 14366 33940 14372 33952
rect 14424 33940 14430 33992
rect 14461 33983 14519 33989
rect 14461 33949 14473 33983
rect 14507 33980 14519 33983
rect 15470 33980 15476 33992
rect 14507 33952 15476 33980
rect 14507 33949 14519 33952
rect 14461 33943 14519 33949
rect 15470 33940 15476 33952
rect 15528 33940 15534 33992
rect 15930 33980 15936 33992
rect 15891 33952 15936 33980
rect 15930 33940 15936 33952
rect 15988 33940 15994 33992
rect 16117 33983 16175 33989
rect 16117 33949 16129 33983
rect 16163 33949 16175 33983
rect 16117 33943 16175 33949
rect 12529 33915 12587 33921
rect 12529 33881 12541 33915
rect 12575 33912 12587 33915
rect 12894 33912 12900 33924
rect 12575 33884 12900 33912
rect 12575 33881 12587 33884
rect 12529 33875 12587 33881
rect 12894 33872 12900 33884
rect 12952 33872 12958 33924
rect 15488 33912 15516 33940
rect 16132 33912 16160 33943
rect 15488 33884 16160 33912
rect 9674 33844 9680 33856
rect 9635 33816 9680 33844
rect 9674 33804 9680 33816
rect 9732 33804 9738 33856
rect 13541 33847 13599 33853
rect 13541 33813 13553 33847
rect 13587 33844 13599 33847
rect 13998 33844 14004 33856
rect 13587 33816 14004 33844
rect 13587 33813 13599 33816
rect 13541 33807 13599 33813
rect 13998 33804 14004 33816
rect 14056 33804 14062 33856
rect 14642 33844 14648 33856
rect 14603 33816 14648 33844
rect 14642 33804 14648 33816
rect 14700 33804 14706 33856
rect 16025 33847 16083 33853
rect 16025 33813 16037 33847
rect 16071 33844 16083 33847
rect 16114 33844 16120 33856
rect 16071 33816 16120 33844
rect 16071 33813 16083 33816
rect 16025 33807 16083 33813
rect 16114 33804 16120 33816
rect 16172 33804 16178 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 15930 33600 15936 33652
rect 15988 33640 15994 33652
rect 16117 33643 16175 33649
rect 16117 33640 16129 33643
rect 15988 33612 16129 33640
rect 15988 33600 15994 33612
rect 16117 33609 16129 33612
rect 16163 33609 16175 33643
rect 16117 33603 16175 33609
rect 9674 33532 9680 33584
rect 9732 33572 9738 33584
rect 9830 33575 9888 33581
rect 9830 33572 9842 33575
rect 9732 33544 9842 33572
rect 9732 33532 9738 33544
rect 9830 33541 9842 33544
rect 9876 33541 9888 33575
rect 9830 33535 9888 33541
rect 7736 33507 7794 33513
rect 7736 33473 7748 33507
rect 7782 33504 7794 33507
rect 8294 33504 8300 33516
rect 7782 33476 8300 33504
rect 7782 33473 7794 33476
rect 7736 33467 7794 33473
rect 8294 33464 8300 33476
rect 8352 33464 8358 33516
rect 12618 33504 12624 33516
rect 12579 33476 12624 33504
rect 12618 33464 12624 33476
rect 12676 33464 12682 33516
rect 13814 33464 13820 33516
rect 13872 33504 13878 33516
rect 14257 33507 14315 33513
rect 14257 33504 14269 33507
rect 13872 33476 14269 33504
rect 13872 33464 13878 33476
rect 14257 33473 14269 33476
rect 14303 33473 14315 33507
rect 14257 33467 14315 33473
rect 15286 33464 15292 33516
rect 15344 33504 15350 33516
rect 15841 33507 15899 33513
rect 15841 33504 15853 33507
rect 15344 33476 15853 33504
rect 15344 33464 15350 33476
rect 15841 33473 15853 33476
rect 15887 33473 15899 33507
rect 15841 33467 15899 33473
rect 7469 33439 7527 33445
rect 7469 33405 7481 33439
rect 7515 33405 7527 33439
rect 9585 33439 9643 33445
rect 9585 33436 9597 33439
rect 7469 33399 7527 33405
rect 8496 33408 9597 33436
rect 7484 33300 7512 33399
rect 8110 33300 8116 33312
rect 7484 33272 8116 33300
rect 8110 33260 8116 33272
rect 8168 33300 8174 33312
rect 8496 33300 8524 33408
rect 9585 33405 9597 33408
rect 9631 33405 9643 33439
rect 9585 33399 9643 33405
rect 12066 33396 12072 33448
rect 12124 33436 12130 33448
rect 12345 33439 12403 33445
rect 12345 33436 12357 33439
rect 12124 33408 12357 33436
rect 12124 33396 12130 33408
rect 12345 33405 12357 33408
rect 12391 33405 12403 33439
rect 13998 33436 14004 33448
rect 13911 33408 14004 33436
rect 12345 33399 12403 33405
rect 13998 33396 14004 33408
rect 14056 33396 14062 33448
rect 16117 33439 16175 33445
rect 16117 33405 16129 33439
rect 16163 33436 16175 33439
rect 16206 33436 16212 33448
rect 16163 33408 16212 33436
rect 16163 33405 16175 33408
rect 16117 33399 16175 33405
rect 16206 33396 16212 33408
rect 16264 33396 16270 33448
rect 8846 33300 8852 33312
rect 8168 33272 8524 33300
rect 8807 33272 8852 33300
rect 8168 33260 8174 33272
rect 8846 33260 8852 33272
rect 8904 33260 8910 33312
rect 10962 33300 10968 33312
rect 10923 33272 10968 33300
rect 10962 33260 10968 33272
rect 11020 33260 11026 33312
rect 12802 33260 12808 33312
rect 12860 33300 12866 33312
rect 13906 33300 13912 33312
rect 12860 33272 13912 33300
rect 12860 33260 12866 33272
rect 13906 33260 13912 33272
rect 13964 33260 13970 33312
rect 14016 33300 14044 33396
rect 15381 33371 15439 33377
rect 15381 33337 15393 33371
rect 15427 33368 15439 33371
rect 17034 33368 17040 33380
rect 15427 33340 17040 33368
rect 15427 33337 15439 33340
rect 15381 33331 15439 33337
rect 17034 33328 17040 33340
rect 17092 33328 17098 33380
rect 14918 33300 14924 33312
rect 14016 33272 14924 33300
rect 14918 33260 14924 33272
rect 14976 33260 14982 33312
rect 15746 33260 15752 33312
rect 15804 33300 15810 33312
rect 15933 33303 15991 33309
rect 15933 33300 15945 33303
rect 15804 33272 15945 33300
rect 15804 33260 15810 33272
rect 15933 33269 15945 33272
rect 15979 33300 15991 33303
rect 16482 33300 16488 33312
rect 15979 33272 16488 33300
rect 15979 33269 15991 33272
rect 15933 33263 15991 33269
rect 16482 33260 16488 33272
rect 16540 33260 16546 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 8573 33099 8631 33105
rect 8573 33065 8585 33099
rect 8619 33096 8631 33099
rect 9858 33096 9864 33108
rect 8619 33068 9864 33096
rect 8619 33065 8631 33068
rect 8573 33059 8631 33065
rect 9858 33056 9864 33068
rect 9916 33056 9922 33108
rect 12802 33096 12808 33108
rect 9968 33068 12808 33096
rect 9968 33028 9996 33068
rect 12802 33056 12808 33068
rect 12860 33056 12866 33108
rect 12894 33056 12900 33108
rect 12952 33096 12958 33108
rect 16666 33096 16672 33108
rect 12952 33068 16672 33096
rect 12952 33056 12958 33068
rect 8220 33000 9996 33028
rect 8220 32969 8248 33000
rect 7285 32963 7343 32969
rect 7285 32929 7297 32963
rect 7331 32960 7343 32963
rect 8205 32963 8263 32969
rect 8205 32960 8217 32963
rect 7331 32932 8217 32960
rect 7331 32929 7343 32932
rect 7285 32923 7343 32929
rect 8205 32929 8217 32932
rect 8251 32929 8263 32963
rect 8205 32923 8263 32929
rect 8846 32920 8852 32972
rect 8904 32960 8910 32972
rect 9125 32963 9183 32969
rect 9125 32960 9137 32963
rect 8904 32932 9137 32960
rect 8904 32920 8910 32932
rect 9125 32929 9137 32932
rect 9171 32929 9183 32963
rect 15562 32960 15568 32972
rect 9125 32923 9183 32929
rect 13372 32932 15568 32960
rect 7466 32892 7472 32904
rect 7427 32864 7472 32892
rect 7466 32852 7472 32864
rect 7524 32852 7530 32904
rect 8386 32892 8392 32904
rect 8347 32864 8392 32892
rect 8386 32852 8392 32864
rect 8444 32852 8450 32904
rect 9398 32892 9404 32904
rect 9359 32864 9404 32892
rect 9398 32852 9404 32864
rect 9456 32852 9462 32904
rect 10873 32895 10931 32901
rect 10873 32861 10885 32895
rect 10919 32892 10931 32895
rect 10962 32892 10968 32904
rect 10919 32864 10968 32892
rect 10919 32861 10931 32864
rect 10873 32855 10931 32861
rect 10962 32852 10968 32864
rect 11020 32852 11026 32904
rect 11054 32852 11060 32904
rect 11112 32892 11118 32904
rect 11149 32895 11207 32901
rect 11149 32892 11161 32895
rect 11112 32864 11161 32892
rect 11112 32852 11118 32864
rect 11149 32861 11161 32864
rect 11195 32861 11207 32895
rect 11149 32855 11207 32861
rect 12161 32895 12219 32901
rect 12161 32861 12173 32895
rect 12207 32892 12219 32895
rect 12894 32892 12900 32904
rect 12207 32864 12900 32892
rect 12207 32861 12219 32864
rect 12161 32855 12219 32861
rect 12894 32852 12900 32864
rect 12952 32852 12958 32904
rect 12428 32827 12486 32833
rect 12428 32793 12440 32827
rect 12474 32824 12486 32827
rect 12710 32824 12716 32836
rect 12474 32796 12716 32824
rect 12474 32793 12486 32796
rect 12428 32787 12486 32793
rect 12710 32784 12716 32796
rect 12768 32784 12774 32836
rect 7650 32756 7656 32768
rect 7611 32728 7656 32756
rect 7650 32716 7656 32728
rect 7708 32716 7714 32768
rect 10318 32716 10324 32768
rect 10376 32756 10382 32768
rect 13372 32756 13400 32932
rect 14366 32852 14372 32904
rect 14424 32892 14430 32904
rect 14844 32901 14872 32932
rect 15562 32920 15568 32932
rect 15620 32920 15626 32972
rect 16040 32969 16068 33068
rect 16666 33056 16672 33068
rect 16724 33056 16730 33108
rect 16025 32963 16083 32969
rect 16025 32929 16037 32963
rect 16071 32929 16083 32963
rect 16025 32923 16083 32929
rect 14737 32895 14795 32901
rect 14737 32892 14749 32895
rect 14424 32864 14749 32892
rect 14424 32852 14430 32864
rect 14737 32861 14749 32864
rect 14783 32861 14795 32895
rect 14737 32855 14795 32861
rect 14829 32895 14887 32901
rect 14829 32861 14841 32895
rect 14875 32861 14887 32895
rect 15470 32892 15476 32904
rect 14829 32855 14887 32861
rect 15212 32864 15476 32892
rect 14553 32827 14611 32833
rect 14553 32793 14565 32827
rect 14599 32824 14611 32827
rect 15212 32824 15240 32864
rect 15470 32852 15476 32864
rect 15528 32852 15534 32904
rect 16114 32852 16120 32904
rect 16172 32892 16178 32904
rect 16281 32895 16339 32901
rect 16281 32892 16293 32895
rect 16172 32864 16293 32892
rect 16172 32852 16178 32864
rect 16281 32861 16293 32864
rect 16327 32861 16339 32895
rect 38286 32892 38292 32904
rect 38247 32864 38292 32892
rect 16281 32855 16339 32861
rect 38286 32852 38292 32864
rect 38344 32852 38350 32904
rect 15378 32824 15384 32836
rect 14599 32796 15240 32824
rect 15291 32796 15384 32824
rect 14599 32793 14611 32796
rect 14553 32787 14611 32793
rect 15378 32784 15384 32796
rect 15436 32824 15442 32836
rect 18046 32824 18052 32836
rect 15436 32796 18052 32824
rect 15436 32784 15442 32796
rect 18046 32784 18052 32796
rect 18104 32784 18110 32836
rect 13538 32756 13544 32768
rect 10376 32728 13400 32756
rect 13499 32728 13544 32756
rect 10376 32716 10382 32728
rect 13538 32716 13544 32728
rect 13596 32716 13602 32768
rect 14826 32756 14832 32768
rect 14787 32728 14832 32756
rect 14826 32716 14832 32728
rect 14884 32716 14890 32768
rect 15470 32716 15476 32768
rect 15528 32756 15534 32768
rect 16022 32756 16028 32768
rect 15528 32728 16028 32756
rect 15528 32716 15534 32728
rect 16022 32716 16028 32728
rect 16080 32716 16086 32768
rect 16758 32716 16764 32768
rect 16816 32756 16822 32768
rect 17405 32759 17463 32765
rect 17405 32756 17417 32759
rect 16816 32728 17417 32756
rect 16816 32716 16822 32728
rect 17405 32725 17417 32728
rect 17451 32725 17463 32759
rect 17405 32719 17463 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 7282 32512 7288 32564
rect 7340 32552 7346 32564
rect 7340 32524 8248 32552
rect 7340 32512 7346 32524
rect 8110 32484 8116 32496
rect 6564 32456 8116 32484
rect 6564 32425 6592 32456
rect 8110 32444 8116 32456
rect 8168 32444 8174 32496
rect 8220 32484 8248 32524
rect 8294 32512 8300 32564
rect 8352 32552 8358 32564
rect 8389 32555 8447 32561
rect 8389 32552 8401 32555
rect 8352 32524 8401 32552
rect 8352 32512 8358 32524
rect 8389 32521 8401 32524
rect 8435 32521 8447 32555
rect 8754 32552 8760 32564
rect 8389 32515 8447 32521
rect 8496 32524 8760 32552
rect 8496 32484 8524 32524
rect 8754 32512 8760 32524
rect 8812 32552 8818 32564
rect 11054 32552 11060 32564
rect 8812 32524 11060 32552
rect 8812 32512 8818 32524
rect 11054 32512 11060 32524
rect 11112 32512 11118 32564
rect 12710 32552 12716 32564
rect 12671 32524 12716 32552
rect 12710 32512 12716 32524
rect 12768 32512 12774 32564
rect 13633 32555 13691 32561
rect 13633 32521 13645 32555
rect 13679 32552 13691 32555
rect 14366 32552 14372 32564
rect 13679 32524 14372 32552
rect 13679 32521 13691 32524
rect 13633 32515 13691 32521
rect 14366 32512 14372 32524
rect 14424 32512 14430 32564
rect 16022 32512 16028 32564
rect 16080 32552 16086 32564
rect 17221 32555 17279 32561
rect 17221 32552 17233 32555
rect 16080 32524 17233 32552
rect 16080 32512 16086 32524
rect 17221 32521 17233 32524
rect 17267 32521 17279 32555
rect 17221 32515 17279 32521
rect 10318 32484 10324 32496
rect 8220 32456 8524 32484
rect 9416 32456 10324 32484
rect 6822 32425 6828 32428
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32385 6607 32419
rect 6816 32416 6828 32425
rect 6783 32388 6828 32416
rect 6549 32379 6607 32385
rect 6816 32379 6828 32388
rect 6822 32376 6828 32379
rect 6880 32376 6886 32428
rect 7650 32376 7656 32428
rect 7708 32416 7714 32428
rect 9416 32425 9444 32456
rect 10318 32444 10324 32456
rect 10376 32444 10382 32496
rect 13449 32487 13507 32493
rect 10428 32456 13400 32484
rect 8573 32419 8631 32425
rect 8573 32416 8585 32419
rect 7708 32388 8585 32416
rect 7708 32376 7714 32388
rect 8573 32385 8585 32388
rect 8619 32385 8631 32419
rect 8573 32379 8631 32385
rect 9401 32419 9459 32425
rect 9401 32385 9413 32419
rect 9447 32385 9459 32419
rect 9401 32379 9459 32385
rect 9490 32376 9496 32428
rect 9548 32416 9554 32428
rect 10428 32425 10456 32456
rect 10229 32419 10287 32425
rect 10229 32416 10241 32419
rect 9548 32388 10241 32416
rect 9548 32376 9554 32388
rect 10229 32385 10241 32388
rect 10275 32385 10287 32419
rect 10229 32379 10287 32385
rect 10413 32419 10471 32425
rect 10413 32385 10425 32419
rect 10459 32385 10471 32419
rect 10413 32379 10471 32385
rect 10873 32419 10931 32425
rect 10873 32385 10885 32419
rect 10919 32385 10931 32419
rect 11054 32416 11060 32428
rect 11015 32388 11060 32416
rect 10873 32379 10931 32385
rect 8846 32308 8852 32360
rect 8904 32348 8910 32360
rect 9309 32351 9367 32357
rect 9309 32348 9321 32351
rect 8904 32320 9321 32348
rect 8904 32308 8910 32320
rect 9309 32317 9321 32320
rect 9355 32317 9367 32351
rect 10888 32348 10916 32379
rect 11054 32376 11060 32388
rect 11112 32376 11118 32428
rect 11885 32419 11943 32425
rect 11885 32385 11897 32419
rect 11931 32416 11943 32419
rect 12710 32416 12716 32428
rect 11931 32388 12716 32416
rect 11931 32385 11943 32388
rect 11885 32379 11943 32385
rect 12710 32376 12716 32388
rect 12768 32376 12774 32428
rect 12897 32419 12955 32425
rect 12897 32385 12909 32419
rect 12943 32416 12955 32419
rect 13170 32416 13176 32428
rect 12943 32388 13176 32416
rect 12943 32385 12955 32388
rect 12897 32379 12955 32385
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 9309 32311 9367 32317
rect 9600 32320 10916 32348
rect 8570 32240 8576 32292
rect 8628 32280 8634 32292
rect 9600 32280 9628 32320
rect 9766 32280 9772 32292
rect 8628 32252 9628 32280
rect 9727 32252 9772 32280
rect 8628 32240 8634 32252
rect 9766 32240 9772 32252
rect 9824 32240 9830 32292
rect 10888 32280 10916 32320
rect 10962 32308 10968 32360
rect 11020 32348 11026 32360
rect 11793 32351 11851 32357
rect 11793 32348 11805 32351
rect 11020 32320 11805 32348
rect 11020 32308 11026 32320
rect 11793 32317 11805 32320
rect 11839 32317 11851 32351
rect 11793 32311 11851 32317
rect 11882 32280 11888 32292
rect 10888 32252 11888 32280
rect 11882 32240 11888 32252
rect 11940 32240 11946 32292
rect 7926 32212 7932 32224
rect 7887 32184 7932 32212
rect 7926 32172 7932 32184
rect 7984 32172 7990 32224
rect 10321 32215 10379 32221
rect 10321 32181 10333 32215
rect 10367 32212 10379 32215
rect 10594 32212 10600 32224
rect 10367 32184 10600 32212
rect 10367 32181 10379 32184
rect 10321 32175 10379 32181
rect 10594 32172 10600 32184
rect 10652 32172 10658 32224
rect 10962 32212 10968 32224
rect 10923 32184 10968 32212
rect 10962 32172 10968 32184
rect 11020 32172 11026 32224
rect 11974 32172 11980 32224
rect 12032 32212 12038 32224
rect 12161 32215 12219 32221
rect 12161 32212 12173 32215
rect 12032 32184 12173 32212
rect 12032 32172 12038 32184
rect 12161 32181 12173 32184
rect 12207 32181 12219 32215
rect 13372 32212 13400 32456
rect 13449 32453 13461 32487
rect 13495 32484 13507 32487
rect 14642 32484 14648 32496
rect 13495 32456 14648 32484
rect 13495 32453 13507 32456
rect 13449 32447 13507 32453
rect 14642 32444 14648 32456
rect 14700 32444 14706 32496
rect 15562 32444 15568 32496
rect 15620 32484 15626 32496
rect 15620 32456 16068 32484
rect 15620 32444 15626 32456
rect 13725 32419 13783 32425
rect 13725 32385 13737 32419
rect 13771 32416 13783 32419
rect 15470 32416 15476 32428
rect 13771 32388 15476 32416
rect 13771 32385 13783 32388
rect 13725 32379 13783 32385
rect 15470 32376 15476 32388
rect 15528 32376 15534 32428
rect 15654 32416 15660 32428
rect 15615 32388 15660 32416
rect 15654 32376 15660 32388
rect 15712 32376 15718 32428
rect 15838 32416 15844 32428
rect 15799 32388 15844 32416
rect 15838 32376 15844 32388
rect 15896 32376 15902 32428
rect 15933 32419 15991 32425
rect 15933 32385 15945 32419
rect 15979 32416 15991 32419
rect 16040 32416 16068 32456
rect 15979 32388 16068 32416
rect 15979 32385 15991 32388
rect 15933 32379 15991 32385
rect 16482 32376 16488 32428
rect 16540 32416 16546 32428
rect 17037 32419 17095 32425
rect 17037 32416 17049 32419
rect 16540 32388 17049 32416
rect 16540 32376 16546 32388
rect 17037 32385 17049 32388
rect 17083 32385 17095 32419
rect 17037 32379 17095 32385
rect 17218 32376 17224 32428
rect 17276 32416 17282 32428
rect 17865 32419 17923 32425
rect 17865 32416 17877 32419
rect 17276 32388 17877 32416
rect 17276 32376 17282 32388
rect 17865 32385 17877 32388
rect 17911 32385 17923 32419
rect 17865 32379 17923 32385
rect 14185 32351 14243 32357
rect 14185 32317 14197 32351
rect 14231 32317 14243 32351
rect 14185 32311 14243 32317
rect 13449 32283 13507 32289
rect 13449 32249 13461 32283
rect 13495 32280 13507 32283
rect 13814 32280 13820 32292
rect 13495 32252 13820 32280
rect 13495 32249 13507 32252
rect 13449 32243 13507 32249
rect 13814 32240 13820 32252
rect 13872 32240 13878 32292
rect 14200 32280 14228 32311
rect 14550 32308 14556 32360
rect 14608 32348 14614 32360
rect 15286 32348 15292 32360
rect 14608 32320 15292 32348
rect 14608 32308 14614 32320
rect 15286 32308 15292 32320
rect 15344 32348 15350 32360
rect 15749 32351 15807 32357
rect 15749 32348 15761 32351
rect 15344 32320 15761 32348
rect 15344 32308 15350 32320
rect 15749 32317 15761 32320
rect 15795 32348 15807 32351
rect 16853 32351 16911 32357
rect 16853 32348 16865 32351
rect 15795 32320 16865 32348
rect 15795 32317 15807 32320
rect 15749 32311 15807 32317
rect 16853 32317 16865 32320
rect 16899 32317 16911 32351
rect 16853 32311 16911 32317
rect 16758 32280 16764 32292
rect 14200 32252 16764 32280
rect 16758 32240 16764 32252
rect 16816 32240 16822 32292
rect 14415 32215 14473 32221
rect 14415 32212 14427 32215
rect 13372 32184 14427 32212
rect 12161 32175 12219 32181
rect 14415 32181 14427 32184
rect 14461 32212 14473 32215
rect 14550 32212 14556 32224
rect 14461 32184 14556 32212
rect 14461 32181 14473 32184
rect 14415 32175 14473 32181
rect 14550 32172 14556 32184
rect 14608 32172 14614 32224
rect 15473 32215 15531 32221
rect 15473 32181 15485 32215
rect 15519 32212 15531 32215
rect 16206 32212 16212 32224
rect 15519 32184 16212 32212
rect 15519 32181 15531 32184
rect 15473 32175 15531 32181
rect 16206 32172 16212 32184
rect 16264 32172 16270 32224
rect 17678 32212 17684 32224
rect 17639 32184 17684 32212
rect 17678 32172 17684 32184
rect 17736 32172 17742 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 8389 32011 8447 32017
rect 8389 31977 8401 32011
rect 8435 32008 8447 32011
rect 8662 32008 8668 32020
rect 8435 31980 8668 32008
rect 8435 31977 8447 31980
rect 8389 31971 8447 31977
rect 8662 31968 8668 31980
rect 8720 32008 8726 32020
rect 9398 32008 9404 32020
rect 8720 31980 9404 32008
rect 8720 31968 8726 31980
rect 9398 31968 9404 31980
rect 9456 31968 9462 32020
rect 9493 32011 9551 32017
rect 9493 31977 9505 32011
rect 9539 31977 9551 32011
rect 12986 32008 12992 32020
rect 12947 31980 12992 32008
rect 9493 31971 9551 31977
rect 5169 31943 5227 31949
rect 5169 31909 5181 31943
rect 5215 31940 5227 31943
rect 6362 31940 6368 31952
rect 5215 31912 6368 31940
rect 5215 31909 5227 31912
rect 5169 31903 5227 31909
rect 6362 31900 6368 31912
rect 6420 31900 6426 31952
rect 6454 31900 6460 31952
rect 6512 31940 6518 31952
rect 7926 31940 7932 31952
rect 6512 31912 7932 31940
rect 6512 31900 6518 31912
rect 7926 31900 7932 31912
rect 7984 31900 7990 31952
rect 8570 31940 8576 31952
rect 8531 31912 8576 31940
rect 8570 31900 8576 31912
rect 8628 31900 8634 31952
rect 9214 31900 9220 31952
rect 9272 31940 9278 31952
rect 9508 31940 9536 31971
rect 12986 31968 12992 31980
rect 13044 31968 13050 32020
rect 13170 32008 13176 32020
rect 13131 31980 13176 32008
rect 13170 31968 13176 31980
rect 13228 31968 13234 32020
rect 14829 32011 14887 32017
rect 14829 31977 14841 32011
rect 14875 32008 14887 32011
rect 27154 32008 27160 32020
rect 14875 31980 27160 32008
rect 14875 31977 14887 31980
rect 14829 31971 14887 31977
rect 27154 31968 27160 31980
rect 27212 31968 27218 32020
rect 9272 31912 9536 31940
rect 9272 31900 9278 31912
rect 14366 31900 14372 31952
rect 14424 31940 14430 31952
rect 15930 31940 15936 31952
rect 14424 31912 15936 31940
rect 14424 31900 14430 31912
rect 5368 31844 6684 31872
rect 2593 31807 2651 31813
rect 2593 31773 2605 31807
rect 2639 31804 2651 31807
rect 2774 31804 2780 31816
rect 2639 31776 2780 31804
rect 2639 31773 2651 31776
rect 2593 31767 2651 31773
rect 2774 31764 2780 31776
rect 2832 31764 2838 31816
rect 2869 31807 2927 31813
rect 2869 31773 2881 31807
rect 2915 31773 2927 31807
rect 5166 31804 5172 31816
rect 5127 31776 5172 31804
rect 2869 31767 2927 31773
rect 2498 31696 2504 31748
rect 2556 31736 2562 31748
rect 2884 31736 2912 31767
rect 5166 31764 5172 31776
rect 5224 31764 5230 31816
rect 5368 31813 5396 31844
rect 6656 31816 6684 31844
rect 9674 31832 9680 31884
rect 9732 31872 9738 31884
rect 9861 31875 9919 31881
rect 9861 31872 9873 31875
rect 9732 31844 9873 31872
rect 9732 31832 9738 31844
rect 9861 31841 9873 31844
rect 9907 31872 9919 31875
rect 10318 31872 10324 31884
rect 9907 31844 10324 31872
rect 9907 31841 9919 31844
rect 9861 31835 9919 31841
rect 10318 31832 10324 31844
rect 10376 31832 10382 31884
rect 10962 31832 10968 31884
rect 11020 31872 11026 31884
rect 11882 31872 11888 31884
rect 11020 31844 11652 31872
rect 11843 31844 11888 31872
rect 11020 31832 11026 31844
rect 5353 31807 5411 31813
rect 5353 31773 5365 31807
rect 5399 31773 5411 31807
rect 5810 31804 5816 31816
rect 5771 31776 5816 31804
rect 5353 31767 5411 31773
rect 5810 31764 5816 31776
rect 5868 31764 5874 31816
rect 5997 31807 6055 31813
rect 5997 31773 6009 31807
rect 6043 31773 6055 31807
rect 6454 31804 6460 31816
rect 6415 31776 6460 31804
rect 5997 31767 6055 31773
rect 2556 31708 2912 31736
rect 2556 31696 2562 31708
rect 5442 31696 5448 31748
rect 5500 31736 5506 31748
rect 6012 31736 6040 31767
rect 6454 31764 6460 31776
rect 6512 31764 6518 31816
rect 6638 31764 6644 31816
rect 6696 31804 6702 31816
rect 6733 31807 6791 31813
rect 6733 31804 6745 31807
rect 6696 31776 6745 31804
rect 6696 31764 6702 31776
rect 6733 31773 6745 31776
rect 6779 31804 6791 31807
rect 8018 31804 8024 31816
rect 6779 31776 8024 31804
rect 6779 31773 6791 31776
rect 6733 31767 6791 31773
rect 8018 31764 8024 31776
rect 8076 31804 8082 31816
rect 9401 31807 9459 31813
rect 9401 31804 9413 31807
rect 8076 31776 9413 31804
rect 8076 31764 8082 31776
rect 8220 31745 8248 31776
rect 9401 31773 9413 31776
rect 9447 31804 9459 31807
rect 9582 31804 9588 31816
rect 9447 31776 9588 31804
rect 9447 31773 9459 31776
rect 9401 31767 9459 31773
rect 9582 31764 9588 31776
rect 9640 31764 9646 31816
rect 10134 31764 10140 31816
rect 10192 31804 10198 31816
rect 10594 31804 10600 31816
rect 10192 31776 10600 31804
rect 10192 31764 10198 31776
rect 10594 31764 10600 31776
rect 10652 31764 10658 31816
rect 10873 31807 10931 31813
rect 10873 31773 10885 31807
rect 10919 31804 10931 31807
rect 11054 31804 11060 31816
rect 10919 31776 11060 31804
rect 10919 31773 10931 31776
rect 10873 31767 10931 31773
rect 11054 31764 11060 31776
rect 11112 31764 11118 31816
rect 11146 31764 11152 31816
rect 11204 31804 11210 31816
rect 11624 31813 11652 31844
rect 11882 31832 11888 31844
rect 11940 31832 11946 31884
rect 12710 31832 12716 31884
rect 12768 31872 12774 31884
rect 14182 31872 14188 31884
rect 12768 31844 14188 31872
rect 12768 31832 12774 31844
rect 14182 31832 14188 31844
rect 14240 31872 14246 31884
rect 15470 31872 15476 31884
rect 14240 31844 14780 31872
rect 15431 31844 15476 31872
rect 14240 31832 14246 31844
rect 11517 31807 11575 31813
rect 11517 31804 11529 31807
rect 11204 31776 11529 31804
rect 11204 31764 11210 31776
rect 11517 31773 11529 31776
rect 11563 31773 11575 31807
rect 11517 31767 11575 31773
rect 11609 31807 11667 31813
rect 11609 31773 11621 31807
rect 11655 31773 11667 31807
rect 11609 31767 11667 31773
rect 14277 31807 14335 31813
rect 14277 31773 14289 31807
rect 14323 31804 14335 31807
rect 14366 31804 14372 31816
rect 14323 31776 14372 31804
rect 14323 31773 14335 31776
rect 14277 31767 14335 31773
rect 14366 31764 14372 31776
rect 14424 31764 14430 31816
rect 14642 31804 14648 31816
rect 14603 31776 14648 31804
rect 14642 31764 14648 31776
rect 14700 31764 14706 31816
rect 14752 31804 14780 31844
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 15580 31881 15608 31912
rect 15930 31900 15936 31912
rect 15988 31900 15994 31952
rect 18046 31940 18052 31952
rect 18007 31912 18052 31940
rect 18046 31900 18052 31912
rect 18104 31900 18110 31952
rect 15566 31875 15624 31881
rect 15566 31841 15578 31875
rect 15612 31841 15624 31875
rect 15566 31835 15624 31841
rect 15654 31832 15660 31884
rect 15712 31872 15718 31884
rect 15712 31844 15757 31872
rect 15712 31832 15718 31844
rect 15838 31832 15844 31884
rect 15896 31872 15902 31884
rect 16669 31875 16727 31881
rect 16669 31872 16681 31875
rect 15896 31844 16681 31872
rect 15896 31832 15902 31844
rect 16669 31841 16681 31844
rect 16715 31841 16727 31875
rect 16669 31835 16727 31841
rect 15749 31807 15807 31813
rect 15749 31804 15761 31807
rect 14752 31776 15761 31804
rect 15488 31748 15516 31776
rect 15749 31773 15761 31776
rect 15795 31773 15807 31807
rect 15749 31767 15807 31773
rect 16936 31807 16994 31813
rect 16936 31773 16948 31807
rect 16982 31804 16994 31807
rect 17678 31804 17684 31816
rect 16982 31776 17684 31804
rect 16982 31773 16994 31776
rect 16936 31767 16994 31773
rect 17678 31764 17684 31776
rect 17736 31764 17742 31816
rect 19978 31804 19984 31816
rect 19939 31776 19984 31804
rect 19978 31764 19984 31776
rect 20036 31764 20042 31816
rect 5500 31708 6040 31736
rect 8205 31739 8263 31745
rect 5500 31696 5506 31708
rect 8205 31705 8217 31739
rect 8251 31705 8263 31739
rect 8205 31699 8263 31705
rect 8294 31696 8300 31748
rect 8352 31736 8358 31748
rect 8405 31739 8463 31745
rect 8405 31736 8417 31739
rect 8352 31708 8417 31736
rect 8352 31696 8358 31708
rect 8405 31705 8417 31708
rect 8451 31705 8463 31739
rect 11238 31736 11244 31748
rect 8405 31699 8463 31705
rect 9692 31708 11244 31736
rect 5902 31668 5908 31680
rect 5863 31640 5908 31668
rect 5902 31628 5908 31640
rect 5960 31628 5966 31680
rect 5994 31628 6000 31680
rect 6052 31668 6058 31680
rect 9692 31668 9720 31708
rect 11238 31696 11244 31708
rect 11296 31696 11302 31748
rect 11974 31736 11980 31748
rect 11887 31708 11980 31736
rect 11974 31696 11980 31708
rect 12032 31696 12038 31748
rect 12805 31739 12863 31745
rect 12805 31705 12817 31739
rect 12851 31736 12863 31739
rect 13722 31736 13728 31748
rect 12851 31708 13728 31736
rect 12851 31705 12863 31708
rect 12805 31699 12863 31705
rect 13722 31696 13728 31708
rect 13780 31696 13786 31748
rect 14458 31736 14464 31748
rect 14419 31708 14464 31736
rect 14458 31696 14464 31708
rect 14516 31696 14522 31748
rect 14550 31696 14556 31748
rect 14608 31736 14614 31748
rect 14608 31708 14653 31736
rect 14608 31696 14614 31708
rect 15470 31696 15476 31748
rect 15528 31696 15534 31748
rect 6052 31640 9720 31668
rect 6052 31628 6058 31640
rect 9950 31628 9956 31680
rect 10008 31668 10014 31680
rect 10505 31671 10563 31677
rect 10505 31668 10517 31671
rect 10008 31640 10517 31668
rect 10008 31628 10014 31640
rect 10505 31637 10517 31640
rect 10551 31637 10563 31671
rect 10686 31668 10692 31680
rect 10647 31640 10692 31668
rect 10505 31631 10563 31637
rect 10686 31628 10692 31640
rect 10744 31628 10750 31680
rect 11330 31668 11336 31680
rect 11291 31640 11336 31668
rect 11330 31628 11336 31640
rect 11388 31628 11394 31680
rect 11514 31628 11520 31680
rect 11572 31668 11578 31680
rect 11992 31668 12020 31696
rect 11572 31640 12020 31668
rect 11572 31628 11578 31640
rect 12434 31628 12440 31680
rect 12492 31668 12498 31680
rect 13005 31671 13063 31677
rect 13005 31668 13017 31671
rect 12492 31640 13017 31668
rect 12492 31628 12498 31640
rect 13005 31637 13017 31640
rect 13051 31637 13063 31671
rect 15286 31668 15292 31680
rect 15247 31640 15292 31668
rect 13005 31631 13063 31637
rect 15286 31628 15292 31640
rect 15344 31628 15350 31680
rect 19797 31671 19855 31677
rect 19797 31637 19809 31671
rect 19843 31668 19855 31671
rect 20070 31668 20076 31680
rect 19843 31640 20076 31668
rect 19843 31637 19855 31640
rect 19797 31631 19855 31637
rect 20070 31628 20076 31640
rect 20128 31628 20134 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 2700 31436 5764 31464
rect 1946 31220 1952 31272
rect 2004 31260 2010 31272
rect 2498 31260 2504 31272
rect 2004 31232 2504 31260
rect 2004 31220 2010 31232
rect 2498 31220 2504 31232
rect 2556 31220 2562 31272
rect 2590 31220 2596 31272
rect 2648 31260 2654 31272
rect 2700 31260 2728 31436
rect 2774 31356 2780 31408
rect 2832 31396 2838 31408
rect 5736 31396 5764 31436
rect 5810 31424 5816 31476
rect 5868 31464 5874 31476
rect 6730 31464 6736 31476
rect 5868 31436 6736 31464
rect 5868 31424 5874 31436
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 8110 31464 8116 31476
rect 6840 31436 8116 31464
rect 6840 31396 6868 31436
rect 8110 31424 8116 31436
rect 8168 31424 8174 31476
rect 10505 31467 10563 31473
rect 10505 31433 10517 31467
rect 10551 31464 10563 31467
rect 10551 31436 12296 31464
rect 10551 31433 10563 31436
rect 10505 31427 10563 31433
rect 9766 31396 9772 31408
rect 2832 31368 5672 31396
rect 5736 31368 6868 31396
rect 7484 31368 8616 31396
rect 2832 31356 2838 31368
rect 3786 31328 3792 31340
rect 3747 31300 3792 31328
rect 3786 31288 3792 31300
rect 3844 31288 3850 31340
rect 4080 31337 4108 31368
rect 4065 31331 4123 31337
rect 4065 31297 4077 31331
rect 4111 31297 4123 31331
rect 4065 31291 4123 31297
rect 4982 31288 4988 31340
rect 5040 31328 5046 31340
rect 5261 31331 5319 31337
rect 5261 31328 5273 31331
rect 5040 31300 5273 31328
rect 5040 31288 5046 31300
rect 5261 31297 5273 31300
rect 5307 31297 5319 31331
rect 5644 31328 5672 31368
rect 5994 31328 6000 31340
rect 5644 31300 6000 31328
rect 5261 31291 5319 31297
rect 5994 31288 6000 31300
rect 6052 31288 6058 31340
rect 6638 31328 6644 31340
rect 6599 31300 6644 31328
rect 6638 31288 6644 31300
rect 6696 31288 6702 31340
rect 6825 31331 6883 31337
rect 6825 31297 6837 31331
rect 6871 31297 6883 31331
rect 7282 31328 7288 31340
rect 7243 31300 7288 31328
rect 6825 31291 6883 31297
rect 2777 31263 2835 31269
rect 2777 31260 2789 31263
rect 2648 31232 2789 31260
rect 2648 31220 2654 31232
rect 2777 31229 2789 31232
rect 2823 31229 2835 31263
rect 2777 31223 2835 31229
rect 5353 31263 5411 31269
rect 5353 31229 5365 31263
rect 5399 31260 5411 31263
rect 6454 31260 6460 31272
rect 5399 31232 6460 31260
rect 5399 31229 5411 31232
rect 5353 31223 5411 31229
rect 6454 31220 6460 31232
rect 6512 31220 6518 31272
rect 6840 31260 6868 31291
rect 7282 31288 7288 31300
rect 7340 31288 7346 31340
rect 7484 31337 7512 31368
rect 7469 31331 7527 31337
rect 7469 31297 7481 31331
rect 7515 31297 7527 31331
rect 7469 31291 7527 31297
rect 8018 31288 8024 31340
rect 8076 31328 8082 31340
rect 8159 31331 8217 31337
rect 8159 31328 8171 31331
rect 8076 31300 8171 31328
rect 8076 31288 8082 31300
rect 8159 31297 8171 31300
rect 8205 31297 8217 31331
rect 8291 31328 8297 31340
rect 8252 31300 8297 31328
rect 8159 31291 8217 31297
rect 8291 31288 8297 31300
rect 8349 31288 8355 31340
rect 8588 31337 8616 31368
rect 9600 31368 9772 31396
rect 8394 31331 8452 31337
rect 8394 31297 8406 31331
rect 8440 31328 8452 31331
rect 8573 31331 8631 31337
rect 8440 31300 8524 31328
rect 8440 31297 8452 31300
rect 8394 31291 8452 31297
rect 6564 31232 6868 31260
rect 8496 31260 8524 31300
rect 8573 31297 8585 31331
rect 8619 31328 8631 31331
rect 8662 31328 8668 31340
rect 8619 31300 8668 31328
rect 8619 31297 8631 31300
rect 8573 31291 8631 31297
rect 8662 31288 8668 31300
rect 8720 31288 8726 31340
rect 9600 31337 9628 31368
rect 9766 31356 9772 31368
rect 9824 31356 9830 31408
rect 10778 31396 10784 31408
rect 10739 31368 10784 31396
rect 10778 31356 10784 31368
rect 10836 31356 10842 31408
rect 10962 31356 10968 31408
rect 11020 31405 11026 31408
rect 11020 31399 11049 31405
rect 11037 31365 11049 31399
rect 11020 31359 11049 31365
rect 11020 31356 11026 31359
rect 11238 31356 11244 31408
rect 11296 31396 11302 31408
rect 12158 31396 12164 31408
rect 11296 31368 12164 31396
rect 11296 31356 11302 31368
rect 12158 31356 12164 31368
rect 12216 31356 12222 31408
rect 9585 31331 9643 31337
rect 9585 31297 9597 31331
rect 9631 31297 9643 31331
rect 9585 31291 9643 31297
rect 9674 31288 9680 31340
rect 9732 31328 9738 31340
rect 9732 31300 9777 31328
rect 9732 31288 9738 31300
rect 9858 31288 9864 31340
rect 9916 31328 9922 31340
rect 9916 31300 9961 31328
rect 9916 31288 9922 31300
rect 10594 31288 10600 31340
rect 10652 31328 10658 31340
rect 10689 31331 10747 31337
rect 10689 31328 10701 31331
rect 10652 31300 10701 31328
rect 10652 31288 10658 31300
rect 10689 31297 10701 31300
rect 10735 31297 10747 31331
rect 10689 31291 10747 31297
rect 10873 31331 10931 31337
rect 10873 31297 10885 31331
rect 10919 31328 10931 31331
rect 11882 31328 11888 31340
rect 10919 31300 11284 31328
rect 11843 31300 11888 31328
rect 10919 31297 10931 31300
rect 10873 31291 10931 31297
rect 11256 31272 11284 31300
rect 11882 31288 11888 31300
rect 11940 31288 11946 31340
rect 12268 31337 12296 31436
rect 12434 31424 12440 31476
rect 12492 31464 12498 31476
rect 22465 31467 22523 31473
rect 12492 31436 12537 31464
rect 12492 31424 12498 31436
rect 22465 31433 22477 31467
rect 22511 31464 22523 31467
rect 23293 31467 23351 31473
rect 23293 31464 23305 31467
rect 22511 31436 23305 31464
rect 22511 31433 22523 31436
rect 22465 31427 22523 31433
rect 23293 31433 23305 31436
rect 23339 31433 23351 31467
rect 23293 31427 23351 31433
rect 13262 31396 13268 31408
rect 13223 31368 13268 31396
rect 13262 31356 13268 31368
rect 13320 31356 13326 31408
rect 20070 31405 20076 31408
rect 20064 31359 20076 31405
rect 20128 31396 20134 31408
rect 24397 31399 24455 31405
rect 20128 31368 20164 31396
rect 20070 31356 20076 31359
rect 20128 31356 20134 31368
rect 24397 31365 24409 31399
rect 24443 31396 24455 31399
rect 25314 31396 25320 31408
rect 24443 31368 25320 31396
rect 24443 31365 24455 31368
rect 24397 31359 24455 31365
rect 25314 31356 25320 31368
rect 25372 31356 25378 31408
rect 12253 31331 12311 31337
rect 12253 31297 12265 31331
rect 12299 31297 12311 31331
rect 13078 31328 13084 31340
rect 13039 31300 13084 31328
rect 12253 31291 12311 31297
rect 13078 31288 13084 31300
rect 13136 31288 13142 31340
rect 13170 31288 13176 31340
rect 13228 31328 13234 31340
rect 13228 31300 13273 31328
rect 13228 31288 13234 31300
rect 14366 31288 14372 31340
rect 14424 31328 14430 31340
rect 15105 31331 15163 31337
rect 15105 31328 15117 31331
rect 14424 31300 15117 31328
rect 14424 31288 14430 31300
rect 15105 31297 15117 31300
rect 15151 31297 15163 31331
rect 16298 31328 16304 31340
rect 16259 31300 16304 31328
rect 15105 31291 15163 31297
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 17310 31328 17316 31340
rect 17271 31300 17316 31328
rect 17310 31288 17316 31300
rect 17368 31288 17374 31340
rect 17862 31288 17868 31340
rect 17920 31328 17926 31340
rect 18213 31331 18271 31337
rect 18213 31328 18225 31331
rect 17920 31300 18225 31328
rect 17920 31288 17926 31300
rect 18213 31297 18225 31300
rect 18259 31297 18271 31331
rect 22002 31328 22008 31340
rect 21963 31300 22008 31328
rect 18213 31291 18271 31297
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 23106 31328 23112 31340
rect 23067 31300 23112 31328
rect 23106 31288 23112 31300
rect 23164 31288 23170 31340
rect 23382 31328 23388 31340
rect 23343 31300 23388 31328
rect 23382 31288 23388 31300
rect 23440 31288 23446 31340
rect 24854 31328 24860 31340
rect 24596 31300 24860 31328
rect 8754 31260 8760 31272
rect 8496 31232 8760 31260
rect 6564 31204 6592 31232
rect 8754 31220 8760 31232
rect 8812 31220 8818 31272
rect 9490 31220 9496 31272
rect 9548 31260 9554 31272
rect 9953 31263 10011 31269
rect 9953 31260 9965 31263
rect 9548 31232 9965 31260
rect 9548 31220 9554 31232
rect 9953 31229 9965 31232
rect 9999 31229 10011 31263
rect 11146 31260 11152 31272
rect 11107 31232 11152 31260
rect 9953 31223 10011 31229
rect 11146 31220 11152 31232
rect 11204 31220 11210 31272
rect 11238 31220 11244 31272
rect 11296 31220 11302 31272
rect 11793 31263 11851 31269
rect 11793 31229 11805 31263
rect 11839 31260 11851 31263
rect 13449 31263 13507 31269
rect 13449 31260 13461 31263
rect 11839 31232 13461 31260
rect 11839 31229 11851 31232
rect 11793 31223 11851 31229
rect 13449 31229 13461 31232
rect 13495 31229 13507 31263
rect 13449 31223 13507 31229
rect 14829 31263 14887 31269
rect 14829 31229 14841 31263
rect 14875 31229 14887 31263
rect 14829 31223 14887 31229
rect 17957 31263 18015 31269
rect 17957 31229 17969 31263
rect 18003 31229 18015 31263
rect 17957 31223 18015 31229
rect 6546 31152 6552 31204
rect 6604 31152 6610 31204
rect 8570 31152 8576 31204
rect 8628 31192 8634 31204
rect 12897 31195 12955 31201
rect 8628 31164 12434 31192
rect 8628 31152 8634 31164
rect 5629 31127 5687 31133
rect 5629 31093 5641 31127
rect 5675 31124 5687 31127
rect 5718 31124 5724 31136
rect 5675 31096 5724 31124
rect 5675 31093 5687 31096
rect 5629 31087 5687 31093
rect 5718 31084 5724 31096
rect 5776 31084 5782 31136
rect 7285 31127 7343 31133
rect 7285 31093 7297 31127
rect 7331 31124 7343 31127
rect 7742 31124 7748 31136
rect 7331 31096 7748 31124
rect 7331 31093 7343 31096
rect 7285 31087 7343 31093
rect 7742 31084 7748 31096
rect 7800 31084 7806 31136
rect 7929 31127 7987 31133
rect 7929 31093 7941 31127
rect 7975 31124 7987 31127
rect 8018 31124 8024 31136
rect 7975 31096 8024 31124
rect 7975 31093 7987 31096
rect 7929 31087 7987 31093
rect 8018 31084 8024 31096
rect 8076 31084 8082 31136
rect 10042 31124 10048 31136
rect 10003 31096 10048 31124
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 12161 31127 12219 31133
rect 12161 31124 12173 31127
rect 11388 31096 12173 31124
rect 11388 31084 11394 31096
rect 12161 31093 12173 31096
rect 12207 31093 12219 31127
rect 12406 31124 12434 31164
rect 12897 31161 12909 31195
rect 12943 31192 12955 31195
rect 13538 31192 13544 31204
rect 12943 31164 13544 31192
rect 12943 31161 12955 31164
rect 12897 31155 12955 31161
rect 13538 31152 13544 31164
rect 13596 31152 13602 31204
rect 14366 31152 14372 31204
rect 14424 31192 14430 31204
rect 14844 31192 14872 31223
rect 14424 31164 14872 31192
rect 17497 31195 17555 31201
rect 14424 31152 14430 31164
rect 17497 31161 17509 31195
rect 17543 31192 17555 31195
rect 17972 31192 18000 31223
rect 18966 31220 18972 31272
rect 19024 31260 19030 31272
rect 24596 31269 24624 31300
rect 24854 31288 24860 31300
rect 24912 31288 24918 31340
rect 19797 31263 19855 31269
rect 19797 31260 19809 31263
rect 19024 31232 19809 31260
rect 19024 31220 19030 31232
rect 19797 31229 19809 31232
rect 19843 31229 19855 31263
rect 19797 31223 19855 31229
rect 24581 31263 24639 31269
rect 24581 31229 24593 31263
rect 24627 31229 24639 31263
rect 24762 31260 24768 31272
rect 24723 31232 24768 31260
rect 24581 31223 24639 31229
rect 24762 31220 24768 31232
rect 24820 31220 24826 31272
rect 23014 31192 23020 31204
rect 17543 31164 18000 31192
rect 17543 31161 17555 31164
rect 17497 31155 17555 31161
rect 14458 31124 14464 31136
rect 12406 31096 14464 31124
rect 12161 31087 12219 31093
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 14826 31084 14832 31136
rect 14884 31124 14890 31136
rect 16022 31124 16028 31136
rect 14884 31096 16028 31124
rect 14884 31084 14890 31096
rect 16022 31084 16028 31096
rect 16080 31084 16086 31136
rect 16117 31127 16175 31133
rect 16117 31093 16129 31127
rect 16163 31124 16175 31127
rect 16942 31124 16948 31136
rect 16163 31096 16948 31124
rect 16163 31093 16175 31096
rect 16117 31087 16175 31093
rect 16942 31084 16948 31096
rect 17000 31084 17006 31136
rect 17972 31124 18000 31164
rect 20732 31164 23020 31192
rect 18874 31124 18880 31136
rect 17972 31096 18880 31124
rect 18874 31084 18880 31096
rect 18932 31084 18938 31136
rect 19337 31127 19395 31133
rect 19337 31093 19349 31127
rect 19383 31124 19395 31127
rect 19426 31124 19432 31136
rect 19383 31096 19432 31124
rect 19383 31093 19395 31096
rect 19337 31087 19395 31093
rect 19426 31084 19432 31096
rect 19484 31124 19490 31136
rect 20732 31124 20760 31164
rect 23014 31152 23020 31164
rect 23072 31152 23078 31204
rect 24397 31195 24455 31201
rect 24397 31161 24409 31195
rect 24443 31192 24455 31195
rect 32950 31192 32956 31204
rect 24443 31164 32956 31192
rect 24443 31161 24455 31164
rect 24397 31155 24455 31161
rect 32950 31152 32956 31164
rect 33008 31152 33014 31204
rect 19484 31096 20760 31124
rect 19484 31084 19490 31096
rect 20898 31084 20904 31136
rect 20956 31124 20962 31136
rect 21177 31127 21235 31133
rect 21177 31124 21189 31127
rect 20956 31096 21189 31124
rect 20956 31084 20962 31096
rect 21177 31093 21189 31096
rect 21223 31124 21235 31127
rect 22002 31124 22008 31136
rect 21223 31096 22008 31124
rect 21223 31093 21235 31096
rect 21177 31087 21235 31093
rect 22002 31084 22008 31096
rect 22060 31084 22066 31136
rect 22278 31124 22284 31136
rect 22239 31096 22284 31124
rect 22278 31084 22284 31096
rect 22336 31084 22342 31136
rect 22925 31127 22983 31133
rect 22925 31093 22937 31127
rect 22971 31124 22983 31127
rect 23198 31124 23204 31136
rect 22971 31096 23204 31124
rect 22971 31093 22983 31096
rect 22925 31087 22983 31093
rect 23198 31084 23204 31096
rect 23256 31084 23262 31136
rect 24670 31084 24676 31136
rect 24728 31124 24734 31136
rect 24728 31096 24773 31124
rect 24728 31084 24734 31096
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 11698 30920 11704 30932
rect 6104 30892 6776 30920
rect 6104 30852 6132 30892
rect 4724 30824 6132 30852
rect 2409 30787 2467 30793
rect 2409 30753 2421 30787
rect 2455 30784 2467 30787
rect 2590 30784 2596 30796
rect 2455 30756 2596 30784
rect 2455 30753 2467 30756
rect 2409 30747 2467 30753
rect 2590 30744 2596 30756
rect 2648 30744 2654 30796
rect 4724 30784 4752 30824
rect 4632 30756 4752 30784
rect 2130 30676 2136 30728
rect 2188 30716 2194 30728
rect 4632 30725 4660 30756
rect 5718 30744 5724 30796
rect 5776 30784 5782 30796
rect 6104 30793 6132 30824
rect 6549 30855 6607 30861
rect 6549 30821 6561 30855
rect 6595 30852 6607 30855
rect 6638 30852 6644 30864
rect 6595 30824 6644 30852
rect 6595 30821 6607 30824
rect 6549 30815 6607 30821
rect 6638 30812 6644 30824
rect 6696 30812 6702 30864
rect 6748 30852 6776 30892
rect 7668 30892 11704 30920
rect 7668 30852 7696 30892
rect 11698 30880 11704 30892
rect 11756 30880 11762 30932
rect 11882 30920 11888 30932
rect 11843 30892 11888 30920
rect 11882 30880 11888 30892
rect 11940 30880 11946 30932
rect 12529 30923 12587 30929
rect 12529 30889 12541 30923
rect 12575 30920 12587 30923
rect 12986 30920 12992 30932
rect 12575 30892 12992 30920
rect 12575 30889 12587 30892
rect 12529 30883 12587 30889
rect 12986 30880 12992 30892
rect 13044 30880 13050 30932
rect 14645 30923 14703 30929
rect 14645 30889 14657 30923
rect 14691 30920 14703 30923
rect 15286 30920 15292 30932
rect 14691 30892 15292 30920
rect 14691 30889 14703 30892
rect 14645 30883 14703 30889
rect 15286 30880 15292 30892
rect 15344 30880 15350 30932
rect 15473 30923 15531 30929
rect 15473 30889 15485 30923
rect 15519 30889 15531 30923
rect 15473 30883 15531 30889
rect 15657 30923 15715 30929
rect 15657 30889 15669 30923
rect 15703 30920 15715 30923
rect 15746 30920 15752 30932
rect 15703 30892 15752 30920
rect 15703 30889 15715 30892
rect 15657 30883 15715 30889
rect 6748 30824 7696 30852
rect 10042 30812 10048 30864
rect 10100 30852 10106 30864
rect 15488 30852 15516 30883
rect 15746 30880 15752 30892
rect 15804 30880 15810 30932
rect 16206 30880 16212 30932
rect 16264 30920 16270 30932
rect 16301 30923 16359 30929
rect 16301 30920 16313 30923
rect 16264 30892 16313 30920
rect 16264 30880 16270 30892
rect 16301 30889 16313 30892
rect 16347 30889 16359 30923
rect 16301 30883 16359 30889
rect 16485 30923 16543 30929
rect 16485 30889 16497 30923
rect 16531 30920 16543 30923
rect 17218 30920 17224 30932
rect 16531 30892 17224 30920
rect 16531 30889 16543 30892
rect 16485 30883 16543 30889
rect 17218 30880 17224 30892
rect 17276 30880 17282 30932
rect 17862 30920 17868 30932
rect 17823 30892 17868 30920
rect 17862 30880 17868 30892
rect 17920 30880 17926 30932
rect 18693 30923 18751 30929
rect 18693 30889 18705 30923
rect 18739 30920 18751 30923
rect 19797 30923 19855 30929
rect 19797 30920 19809 30923
rect 18739 30892 19809 30920
rect 18739 30889 18751 30892
rect 18693 30883 18751 30889
rect 19797 30889 19809 30892
rect 19843 30889 19855 30923
rect 19797 30883 19855 30889
rect 24581 30923 24639 30929
rect 24581 30889 24593 30923
rect 24627 30920 24639 30923
rect 24670 30920 24676 30932
rect 24627 30892 24676 30920
rect 24627 30889 24639 30892
rect 24581 30883 24639 30889
rect 24670 30880 24676 30892
rect 24728 30880 24734 30932
rect 15838 30852 15844 30864
rect 10100 30824 11192 30852
rect 15488 30824 15844 30852
rect 10100 30812 10106 30824
rect 5905 30787 5963 30793
rect 5905 30784 5917 30787
rect 5776 30756 5917 30784
rect 5776 30744 5782 30756
rect 5905 30753 5917 30756
rect 5951 30753 5963 30787
rect 5905 30747 5963 30753
rect 6089 30787 6147 30793
rect 6089 30753 6101 30787
rect 6135 30753 6147 30787
rect 6089 30747 6147 30753
rect 2685 30719 2743 30725
rect 2685 30716 2697 30719
rect 2188 30688 2697 30716
rect 2188 30676 2194 30688
rect 2685 30685 2697 30688
rect 2731 30685 2743 30719
rect 2685 30679 2743 30685
rect 4617 30719 4675 30725
rect 4617 30685 4629 30719
rect 4663 30685 4675 30719
rect 4798 30716 4804 30728
rect 4759 30688 4804 30716
rect 4617 30679 4675 30685
rect 4798 30676 4804 30688
rect 4856 30676 4862 30728
rect 4893 30719 4951 30725
rect 4893 30685 4905 30719
rect 4939 30716 4951 30719
rect 5442 30716 5448 30728
rect 4939 30688 5448 30716
rect 4939 30685 4951 30688
rect 4893 30679 4951 30685
rect 5442 30676 5448 30688
rect 5500 30676 5506 30728
rect 5813 30719 5871 30725
rect 5813 30685 5825 30719
rect 5859 30685 5871 30719
rect 5920 30716 5948 30747
rect 6730 30744 6736 30796
rect 6788 30784 6794 30796
rect 6788 30756 7880 30784
rect 6788 30744 6794 30756
rect 6825 30719 6883 30725
rect 6825 30716 6837 30719
rect 5920 30688 6837 30716
rect 5813 30679 5871 30685
rect 6825 30685 6837 30688
rect 6871 30685 6883 30719
rect 7742 30716 7748 30728
rect 7703 30688 7748 30716
rect 6825 30679 6883 30685
rect 5828 30592 5856 30679
rect 7742 30676 7748 30688
rect 7800 30676 7806 30728
rect 7852 30725 7880 30756
rect 8294 30744 8300 30796
rect 8352 30784 8358 30796
rect 8478 30784 8484 30796
rect 8352 30756 8484 30784
rect 8352 30744 8358 30756
rect 8478 30744 8484 30756
rect 8536 30784 8542 30796
rect 9490 30784 9496 30796
rect 8536 30756 9496 30784
rect 8536 30744 8542 30756
rect 9490 30744 9496 30756
rect 9548 30784 9554 30796
rect 9548 30756 9720 30784
rect 9548 30744 9554 30756
rect 7837 30719 7895 30725
rect 7837 30685 7849 30719
rect 7883 30685 7895 30719
rect 8018 30716 8024 30728
rect 7979 30688 8024 30716
rect 7837 30679 7895 30685
rect 8018 30676 8024 30688
rect 8076 30676 8082 30728
rect 8113 30719 8171 30725
rect 8113 30685 8125 30719
rect 8159 30685 8171 30719
rect 9401 30719 9459 30725
rect 9401 30716 9413 30719
rect 8113 30679 8171 30685
rect 9140 30688 9413 30716
rect 6089 30651 6147 30657
rect 6089 30617 6101 30651
rect 6135 30648 6147 30651
rect 6549 30651 6607 30657
rect 6549 30648 6561 30651
rect 6135 30620 6561 30648
rect 6135 30617 6147 30620
rect 6089 30611 6147 30617
rect 6549 30617 6561 30620
rect 6595 30617 6607 30651
rect 6549 30611 6607 30617
rect 7374 30608 7380 30660
rect 7432 30648 7438 30660
rect 8128 30648 8156 30679
rect 7432 30620 8156 30648
rect 7432 30608 7438 30620
rect 4430 30580 4436 30592
rect 4391 30552 4436 30580
rect 4430 30540 4436 30552
rect 4488 30540 4494 30592
rect 5810 30580 5816 30592
rect 5723 30552 5816 30580
rect 5810 30540 5816 30552
rect 5868 30580 5874 30592
rect 6733 30583 6791 30589
rect 6733 30580 6745 30583
rect 5868 30552 6745 30580
rect 5868 30540 5874 30552
rect 6733 30549 6745 30552
rect 6779 30549 6791 30583
rect 6733 30543 6791 30549
rect 7561 30583 7619 30589
rect 7561 30549 7573 30583
rect 7607 30580 7619 30583
rect 8570 30580 8576 30592
rect 7607 30552 8576 30580
rect 7607 30549 7619 30552
rect 7561 30543 7619 30549
rect 8570 30540 8576 30552
rect 8628 30540 8634 30592
rect 9140 30580 9168 30688
rect 9401 30685 9413 30688
rect 9447 30685 9459 30719
rect 9582 30716 9588 30728
rect 9543 30688 9588 30716
rect 9401 30679 9459 30685
rect 9582 30676 9588 30688
rect 9640 30676 9646 30728
rect 9692 30725 9720 30756
rect 9950 30744 9956 30796
rect 10008 30784 10014 30796
rect 10594 30784 10600 30796
rect 10008 30756 10456 30784
rect 10555 30756 10600 30784
rect 10008 30744 10014 30756
rect 9677 30719 9735 30725
rect 9677 30685 9689 30719
rect 9723 30685 9735 30719
rect 9677 30679 9735 30685
rect 10134 30676 10140 30728
rect 10192 30725 10198 30728
rect 10192 30719 10251 30725
rect 10192 30685 10205 30719
rect 10239 30685 10251 30719
rect 10318 30716 10324 30728
rect 10279 30688 10324 30716
rect 10192 30679 10251 30685
rect 10192 30676 10198 30679
rect 10318 30676 10324 30688
rect 10376 30676 10382 30728
rect 10428 30719 10456 30756
rect 10594 30744 10600 30756
rect 10652 30744 10658 30796
rect 11164 30725 11192 30824
rect 15838 30812 15844 30824
rect 15896 30812 15902 30864
rect 18877 30855 18935 30861
rect 18877 30821 18889 30855
rect 18923 30852 18935 30855
rect 19978 30852 19984 30864
rect 18923 30824 19984 30852
rect 18923 30821 18935 30824
rect 18877 30815 18935 30821
rect 19978 30812 19984 30824
rect 20036 30812 20042 30864
rect 23477 30855 23535 30861
rect 23477 30821 23489 30855
rect 23523 30852 23535 30855
rect 24949 30855 25007 30861
rect 24949 30852 24961 30855
rect 23523 30824 24961 30852
rect 23523 30821 23535 30824
rect 23477 30815 23535 30821
rect 24949 30821 24961 30824
rect 24995 30821 25007 30855
rect 24949 30815 25007 30821
rect 11422 30784 11428 30796
rect 11383 30756 11428 30784
rect 11422 30744 11428 30756
rect 11480 30744 11486 30796
rect 11606 30744 11612 30796
rect 11664 30784 11670 30796
rect 12710 30784 12716 30796
rect 11664 30756 12716 30784
rect 11664 30744 11670 30756
rect 12710 30744 12716 30756
rect 12768 30784 12774 30796
rect 13446 30784 13452 30796
rect 12768 30756 13452 30784
rect 12768 30744 12774 30756
rect 13446 30744 13452 30756
rect 13504 30744 13510 30796
rect 14366 30744 14372 30796
rect 14424 30784 14430 30796
rect 17221 30787 17279 30793
rect 17221 30784 17233 30787
rect 14424 30756 17233 30784
rect 14424 30744 14430 30756
rect 17221 30753 17233 30756
rect 17267 30753 17279 30787
rect 20898 30784 20904 30796
rect 20859 30756 20904 30784
rect 17221 30747 17279 30753
rect 20898 30744 20904 30756
rect 20956 30744 20962 30796
rect 21174 30784 21180 30796
rect 21008 30756 21180 30784
rect 11149 30719 11207 30725
rect 10413 30713 10471 30719
rect 10413 30679 10425 30713
rect 10459 30679 10471 30713
rect 11149 30685 11161 30719
rect 11195 30685 11207 30719
rect 11149 30679 11207 30685
rect 11333 30719 11391 30725
rect 11333 30685 11345 30719
rect 11379 30685 11391 30719
rect 11333 30679 11391 30685
rect 10413 30673 10471 30679
rect 9217 30651 9275 30657
rect 9217 30617 9229 30651
rect 9263 30648 9275 30651
rect 9858 30648 9864 30660
rect 9263 30620 9864 30648
rect 9263 30617 9275 30620
rect 9217 30611 9275 30617
rect 9858 30608 9864 30620
rect 9916 30608 9922 30660
rect 9766 30580 9772 30592
rect 9140 30552 9772 30580
rect 9766 30540 9772 30552
rect 9824 30580 9830 30592
rect 10594 30580 10600 30592
rect 9824 30552 10600 30580
rect 9824 30540 9830 30552
rect 10594 30540 10600 30552
rect 10652 30540 10658 30592
rect 11054 30540 11060 30592
rect 11112 30580 11118 30592
rect 11348 30580 11376 30679
rect 11514 30676 11520 30728
rect 11572 30716 11578 30728
rect 11701 30719 11759 30725
rect 11572 30688 11617 30716
rect 11572 30676 11578 30688
rect 11701 30685 11713 30719
rect 11747 30716 11759 30719
rect 11790 30716 11796 30728
rect 11747 30688 11796 30716
rect 11747 30685 11759 30688
rect 11701 30679 11759 30685
rect 11790 30676 11796 30688
rect 11848 30676 11854 30728
rect 12805 30719 12863 30725
rect 12805 30685 12817 30719
rect 12851 30716 12863 30719
rect 12986 30716 12992 30728
rect 12851 30688 12992 30716
rect 12851 30685 12863 30688
rect 12805 30679 12863 30685
rect 12986 30676 12992 30688
rect 13044 30676 13050 30728
rect 13170 30716 13176 30728
rect 13131 30688 13176 30716
rect 13170 30676 13176 30688
rect 13228 30676 13234 30728
rect 15520 30660 15691 30682
rect 16022 30676 16028 30728
rect 16080 30716 16086 30728
rect 17034 30716 17040 30728
rect 16080 30691 16360 30716
rect 16080 30688 16405 30691
rect 16995 30688 17040 30716
rect 16080 30676 16086 30688
rect 16332 30685 16405 30688
rect 13722 30608 13728 30660
rect 13780 30648 13786 30660
rect 14461 30651 14519 30657
rect 14461 30648 14473 30651
rect 13780 30620 14473 30648
rect 13780 30608 13786 30620
rect 14461 30617 14473 30620
rect 14507 30648 14519 30651
rect 14507 30620 15240 30648
rect 14507 30617 14519 30620
rect 14461 30611 14519 30617
rect 12851 30583 12909 30589
rect 12851 30580 12863 30583
rect 11112 30552 12863 30580
rect 11112 30540 11118 30552
rect 12851 30549 12863 30552
rect 12897 30549 12909 30583
rect 13078 30580 13084 30592
rect 13039 30552 13084 30580
rect 12851 30543 12909 30549
rect 13078 30540 13084 30552
rect 13136 30540 13142 30592
rect 14642 30540 14648 30592
rect 14700 30589 14706 30592
rect 14700 30583 14719 30589
rect 14707 30549 14719 30583
rect 14826 30580 14832 30592
rect 14787 30552 14832 30580
rect 14700 30543 14719 30549
rect 14700 30540 14706 30543
rect 14826 30540 14832 30552
rect 14884 30540 14890 30592
rect 15212 30580 15240 30620
rect 15286 30608 15292 30660
rect 15344 30648 15350 30660
rect 15520 30657 15651 30660
rect 15499 30654 15651 30657
rect 15499 30651 15557 30654
rect 15344 30620 15389 30648
rect 15344 30608 15350 30620
rect 15499 30617 15511 30651
rect 15545 30617 15557 30651
rect 15499 30611 15557 30617
rect 15645 30608 15651 30654
rect 15703 30608 15709 30660
rect 16117 30651 16175 30657
rect 16332 30654 16359 30685
rect 16117 30617 16129 30651
rect 16163 30617 16175 30651
rect 16347 30651 16359 30654
rect 16393 30651 16405 30685
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 18049 30719 18107 30725
rect 18049 30685 18061 30719
rect 18095 30716 18107 30719
rect 18414 30716 18420 30728
rect 18095 30688 18420 30716
rect 18095 30685 18107 30688
rect 18049 30679 18107 30685
rect 18414 30676 18420 30688
rect 18472 30676 18478 30728
rect 20438 30716 20444 30728
rect 20399 30688 20444 30716
rect 20438 30676 20444 30688
rect 20496 30676 20502 30728
rect 16347 30645 16405 30651
rect 18509 30651 18567 30657
rect 16117 30611 16175 30617
rect 18509 30617 18521 30651
rect 18555 30648 18567 30651
rect 19242 30648 19248 30660
rect 18555 30620 19248 30648
rect 18555 30617 18567 30620
rect 18509 30611 18567 30617
rect 16132 30580 16160 30611
rect 18524 30580 18552 30611
rect 19242 30608 19248 30620
rect 19300 30608 19306 30660
rect 19334 30608 19340 30660
rect 19392 30648 19398 30660
rect 19429 30651 19487 30657
rect 19429 30648 19441 30651
rect 19392 30620 19441 30648
rect 19392 30608 19398 30620
rect 19429 30617 19441 30620
rect 19475 30617 19487 30651
rect 19429 30611 19487 30617
rect 19613 30651 19671 30657
rect 19613 30617 19625 30651
rect 19659 30648 19671 30651
rect 21008 30648 21036 30756
rect 21174 30744 21180 30756
rect 21232 30744 21238 30796
rect 23014 30784 23020 30796
rect 22975 30756 23020 30784
rect 23014 30744 23020 30756
rect 23072 30744 23078 30796
rect 22554 30676 22560 30728
rect 22612 30716 22618 30728
rect 23109 30719 23167 30725
rect 23109 30716 23121 30719
rect 22612 30688 23121 30716
rect 22612 30676 22618 30688
rect 23109 30685 23121 30688
rect 23155 30685 23167 30719
rect 23109 30679 23167 30685
rect 24670 30676 24676 30728
rect 24728 30716 24734 30728
rect 24765 30719 24823 30725
rect 24765 30716 24777 30719
rect 24728 30688 24777 30716
rect 24728 30676 24734 30688
rect 24765 30685 24777 30688
rect 24811 30685 24823 30719
rect 25038 30716 25044 30728
rect 24999 30688 25044 30716
rect 24765 30679 24823 30685
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 19659 30620 21036 30648
rect 19659 30617 19671 30620
rect 19613 30611 19671 30617
rect 15212 30552 18552 30580
rect 18690 30540 18696 30592
rect 18748 30589 18754 30592
rect 18748 30583 18767 30589
rect 18755 30549 18767 30583
rect 18748 30543 18767 30549
rect 18748 30540 18754 30543
rect 19058 30540 19064 30592
rect 19116 30580 19122 30592
rect 19628 30580 19656 30611
rect 19116 30552 19656 30580
rect 20257 30583 20315 30589
rect 19116 30540 19122 30552
rect 20257 30549 20269 30583
rect 20303 30580 20315 30583
rect 20346 30580 20352 30592
rect 20303 30552 20352 30580
rect 20303 30549 20315 30552
rect 20257 30543 20315 30549
rect 20346 30540 20352 30552
rect 20404 30540 20410 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 3789 30379 3847 30385
rect 3789 30345 3801 30379
rect 3835 30345 3847 30379
rect 4430 30376 4436 30388
rect 4391 30348 4436 30376
rect 3789 30339 3847 30345
rect 3804 30308 3832 30339
rect 4430 30336 4436 30348
rect 4488 30336 4494 30388
rect 5810 30376 5816 30388
rect 5771 30348 5816 30376
rect 5810 30336 5816 30348
rect 5868 30336 5874 30388
rect 6546 30336 6552 30388
rect 6604 30376 6610 30388
rect 8478 30376 8484 30388
rect 6604 30348 6960 30376
rect 8439 30348 8484 30376
rect 6604 30336 6610 30348
rect 4614 30308 4620 30320
rect 3804 30280 4620 30308
rect 4614 30268 4620 30280
rect 4672 30308 4678 30320
rect 6564 30308 6592 30336
rect 6822 30308 6828 30320
rect 4672 30280 6592 30308
rect 6783 30280 6828 30308
rect 4672 30268 4678 30280
rect 6822 30268 6828 30280
rect 6880 30268 6886 30320
rect 6932 30308 6960 30348
rect 8478 30336 8484 30348
rect 8536 30336 8542 30388
rect 9677 30379 9735 30385
rect 9677 30345 9689 30379
rect 9723 30376 9735 30379
rect 9950 30376 9956 30388
rect 9723 30348 9956 30376
rect 9723 30345 9735 30348
rect 9677 30339 9735 30345
rect 9950 30336 9956 30348
rect 10008 30336 10014 30388
rect 10505 30379 10563 30385
rect 10505 30345 10517 30379
rect 10551 30376 10563 30379
rect 10686 30376 10692 30388
rect 10551 30348 10692 30376
rect 10551 30345 10563 30348
rect 10505 30339 10563 30345
rect 10686 30336 10692 30348
rect 10744 30336 10750 30388
rect 12897 30379 12955 30385
rect 12897 30345 12909 30379
rect 12943 30376 12955 30379
rect 13170 30376 13176 30388
rect 12943 30348 13176 30376
rect 12943 30345 12955 30348
rect 12897 30339 12955 30345
rect 13170 30336 13176 30348
rect 13228 30336 13234 30388
rect 16298 30376 16304 30388
rect 16259 30348 16304 30376
rect 16298 30336 16304 30348
rect 16356 30336 16362 30388
rect 18690 30336 18696 30388
rect 18748 30376 18754 30388
rect 18969 30379 19027 30385
rect 18969 30376 18981 30379
rect 18748 30348 18981 30376
rect 18748 30336 18754 30348
rect 18969 30345 18981 30348
rect 19015 30345 19027 30379
rect 18969 30339 19027 30345
rect 22465 30379 22523 30385
rect 22465 30345 22477 30379
rect 22511 30376 22523 30379
rect 23106 30376 23112 30388
rect 22511 30348 23112 30376
rect 22511 30345 22523 30348
rect 22465 30339 22523 30345
rect 23106 30336 23112 30348
rect 23164 30336 23170 30388
rect 23753 30379 23811 30385
rect 23753 30345 23765 30379
rect 23799 30376 23811 30379
rect 24670 30376 24676 30388
rect 23799 30348 24676 30376
rect 23799 30345 23811 30348
rect 23753 30339 23811 30345
rect 24670 30336 24676 30348
rect 24728 30336 24734 30388
rect 6932 30280 7512 30308
rect 2682 30249 2688 30252
rect 2676 30203 2688 30249
rect 2740 30240 2746 30252
rect 2740 30212 2776 30240
rect 2682 30200 2688 30203
rect 2740 30200 2746 30212
rect 4062 30200 4068 30252
rect 4120 30240 4126 30252
rect 4374 30243 4432 30249
rect 4374 30240 4386 30243
rect 4120 30212 4386 30240
rect 4120 30200 4126 30212
rect 4374 30209 4386 30212
rect 4420 30240 4432 30243
rect 5537 30243 5595 30249
rect 4420 30212 5028 30240
rect 4420 30209 4432 30212
rect 4374 30203 4432 30209
rect 2130 30132 2136 30184
rect 2188 30172 2194 30184
rect 2409 30175 2467 30181
rect 2409 30172 2421 30175
rect 2188 30144 2421 30172
rect 2188 30132 2194 30144
rect 2409 30141 2421 30144
rect 2455 30141 2467 30175
rect 2409 30135 2467 30141
rect 4893 30175 4951 30181
rect 4893 30141 4905 30175
rect 4939 30141 4951 30175
rect 5000 30172 5028 30212
rect 5537 30209 5549 30243
rect 5583 30240 5595 30243
rect 5583 30212 6316 30240
rect 5583 30209 5595 30212
rect 5537 30203 5595 30209
rect 5813 30175 5871 30181
rect 5813 30172 5825 30175
rect 5000 30144 5825 30172
rect 4893 30135 4951 30141
rect 5813 30141 5825 30144
rect 5859 30141 5871 30175
rect 6288 30172 6316 30212
rect 6362 30200 6368 30252
rect 6420 30240 6426 30252
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 6420 30212 6561 30240
rect 6420 30200 6426 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6549 30203 6607 30209
rect 6638 30200 6644 30252
rect 6696 30240 6702 30252
rect 7484 30249 7512 30280
rect 7558 30268 7564 30320
rect 7616 30308 7622 30320
rect 9398 30308 9404 30320
rect 7616 30280 9404 30308
rect 7616 30268 7622 30280
rect 9398 30268 9404 30280
rect 9456 30268 9462 30320
rect 11514 30268 11520 30320
rect 11572 30308 11578 30320
rect 12621 30311 12679 30317
rect 12621 30308 12633 30311
rect 11572 30280 12633 30308
rect 11572 30268 11578 30280
rect 12621 30277 12633 30280
rect 12667 30277 12679 30311
rect 14182 30308 14188 30320
rect 14143 30280 14188 30308
rect 12621 30271 12679 30277
rect 14182 30268 14188 30280
rect 14240 30268 14246 30320
rect 14550 30308 14556 30320
rect 14511 30280 14556 30308
rect 14550 30268 14556 30280
rect 14608 30268 14614 30320
rect 16022 30268 16028 30320
rect 16080 30308 16086 30320
rect 16117 30311 16175 30317
rect 16117 30308 16129 30311
rect 16080 30280 16129 30308
rect 16080 30268 16086 30280
rect 16117 30277 16129 30280
rect 16163 30277 16175 30311
rect 16117 30271 16175 30277
rect 17310 30268 17316 30320
rect 17368 30308 17374 30320
rect 22002 30308 22008 30320
rect 17368 30280 20116 30308
rect 21963 30280 22008 30308
rect 17368 30268 17374 30280
rect 7469 30243 7527 30249
rect 6696 30212 6741 30240
rect 6696 30200 6702 30212
rect 7469 30209 7481 30243
rect 7515 30240 7527 30243
rect 8297 30243 8355 30249
rect 8297 30240 8309 30243
rect 7515 30212 8309 30240
rect 7515 30209 7527 30212
rect 7469 30203 7527 30209
rect 8297 30209 8309 30212
rect 8343 30209 8355 30243
rect 9214 30240 9220 30252
rect 9175 30212 9220 30240
rect 8297 30203 8355 30209
rect 6730 30172 6736 30184
rect 6288 30144 6736 30172
rect 5813 30135 5871 30141
rect 4908 30104 4936 30135
rect 6730 30132 6736 30144
rect 6788 30132 6794 30184
rect 6822 30132 6828 30184
rect 6880 30172 6886 30184
rect 6880 30144 6925 30172
rect 6880 30132 6886 30144
rect 8018 30132 8024 30184
rect 8076 30172 8082 30184
rect 8113 30175 8171 30181
rect 8113 30172 8125 30175
rect 8076 30144 8125 30172
rect 8076 30132 8082 30144
rect 8113 30141 8125 30144
rect 8159 30141 8171 30175
rect 8312 30172 8340 30203
rect 9214 30200 9220 30212
rect 9272 30200 9278 30252
rect 10321 30243 10379 30249
rect 10321 30209 10333 30243
rect 10367 30209 10379 30243
rect 10321 30203 10379 30209
rect 10505 30243 10563 30249
rect 10505 30209 10517 30243
rect 10551 30209 10563 30243
rect 10505 30203 10563 30209
rect 10965 30243 11023 30249
rect 10965 30209 10977 30243
rect 11011 30240 11023 30243
rect 11606 30240 11612 30252
rect 11011 30212 11612 30240
rect 11011 30209 11023 30212
rect 10965 30203 11023 30209
rect 10336 30172 10364 30203
rect 8312 30144 10364 30172
rect 8113 30135 8171 30141
rect 5629 30107 5687 30113
rect 5629 30104 5641 30107
rect 4908 30076 5641 30104
rect 5629 30073 5641 30076
rect 5675 30104 5687 30107
rect 7558 30104 7564 30116
rect 5675 30076 7564 30104
rect 5675 30073 5687 30076
rect 5629 30067 5687 30073
rect 7558 30064 7564 30076
rect 7616 30064 7622 30116
rect 10520 30104 10548 30203
rect 11606 30200 11612 30212
rect 11664 30200 11670 30252
rect 12738 30243 12796 30249
rect 12738 30240 12750 30243
rect 11716 30212 12750 30240
rect 10594 30132 10600 30184
rect 10652 30172 10658 30184
rect 11716 30172 11744 30212
rect 12738 30209 12750 30212
rect 12784 30209 12796 30243
rect 13538 30240 13544 30252
rect 13451 30212 13544 30240
rect 12738 30203 12796 30209
rect 13538 30200 13544 30212
rect 13596 30240 13602 30252
rect 14369 30243 14427 30249
rect 13596 30212 14320 30240
rect 13596 30200 13602 30212
rect 12250 30172 12256 30184
rect 10652 30144 11744 30172
rect 12211 30144 12256 30172
rect 10652 30132 10658 30144
rect 12250 30132 12256 30144
rect 12308 30132 12314 30184
rect 12526 30172 12532 30184
rect 12487 30144 12532 30172
rect 12526 30132 12532 30144
rect 12584 30132 12590 30184
rect 12986 30132 12992 30184
rect 13044 30172 13050 30184
rect 13630 30172 13636 30184
rect 13044 30144 13636 30172
rect 13044 30132 13050 30144
rect 13630 30132 13636 30144
rect 13688 30172 13694 30184
rect 13725 30175 13783 30181
rect 13725 30172 13737 30175
rect 13688 30144 13737 30172
rect 13688 30132 13694 30144
rect 13725 30141 13737 30144
rect 13771 30141 13783 30175
rect 13725 30135 13783 30141
rect 13538 30104 13544 30116
rect 7852 30076 10456 30104
rect 10520 30076 13544 30104
rect 3878 29996 3884 30048
rect 3936 30036 3942 30048
rect 4249 30039 4307 30045
rect 4249 30036 4261 30039
rect 3936 30008 4261 30036
rect 3936 29996 3942 30008
rect 4249 30005 4261 30008
rect 4295 30005 4307 30039
rect 4249 29999 4307 30005
rect 4801 30039 4859 30045
rect 4801 30005 4813 30039
rect 4847 30036 4859 30039
rect 5166 30036 5172 30048
rect 4847 30008 5172 30036
rect 4847 30005 4859 30008
rect 4801 29999 4859 30005
rect 5166 29996 5172 30008
rect 5224 30036 5230 30048
rect 5810 30036 5816 30048
rect 5224 30008 5816 30036
rect 5224 29996 5230 30008
rect 5810 29996 5816 30008
rect 5868 29996 5874 30048
rect 6638 29996 6644 30048
rect 6696 30036 6702 30048
rect 6822 30036 6828 30048
rect 6696 30008 6828 30036
rect 6696 29996 6702 30008
rect 6822 29996 6828 30008
rect 6880 30036 6886 30048
rect 7852 30036 7880 30076
rect 6880 30008 7880 30036
rect 6880 29996 6886 30008
rect 7926 29996 7932 30048
rect 7984 30036 7990 30048
rect 9309 30039 9367 30045
rect 9309 30036 9321 30039
rect 7984 30008 9321 30036
rect 7984 29996 7990 30008
rect 9309 30005 9321 30008
rect 9355 30005 9367 30039
rect 10428 30036 10456 30076
rect 13538 30064 13544 30076
rect 13596 30064 13602 30116
rect 14292 30104 14320 30212
rect 14369 30209 14381 30243
rect 14415 30209 14427 30243
rect 14369 30203 14427 30209
rect 14384 30172 14412 30203
rect 14458 30200 14464 30252
rect 14516 30240 14522 30252
rect 15746 30240 15752 30252
rect 14516 30212 14561 30240
rect 15707 30212 15752 30240
rect 14516 30200 14522 30212
rect 15746 30200 15752 30212
rect 15804 30200 15810 30252
rect 16666 30200 16672 30252
rect 16724 30240 16730 30252
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 16724 30212 16865 30240
rect 16724 30200 16730 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 16853 30203 16911 30209
rect 16942 30200 16948 30252
rect 17000 30240 17006 30252
rect 17109 30243 17167 30249
rect 17109 30240 17121 30243
rect 17000 30212 17121 30240
rect 17000 30200 17006 30212
rect 17109 30209 17121 30212
rect 17155 30209 17167 30243
rect 17109 30203 17167 30209
rect 18877 30243 18935 30249
rect 18877 30209 18889 30243
rect 18923 30209 18935 30243
rect 19058 30240 19064 30252
rect 19019 30212 19064 30240
rect 18877 30203 18935 30209
rect 15102 30172 15108 30184
rect 14384 30144 15108 30172
rect 15102 30132 15108 30144
rect 15160 30172 15166 30184
rect 15562 30172 15568 30184
rect 15160 30144 15568 30172
rect 15160 30132 15166 30144
rect 15562 30132 15568 30144
rect 15620 30132 15626 30184
rect 18892 30172 18920 30203
rect 19058 30200 19064 30212
rect 19116 30200 19122 30252
rect 20088 30249 20116 30280
rect 22002 30268 22008 30280
rect 22060 30268 22066 30320
rect 25314 30308 25320 30320
rect 25275 30280 25320 30308
rect 25314 30268 25320 30280
rect 25372 30268 25378 30320
rect 20346 30249 20352 30252
rect 20073 30243 20131 30249
rect 20073 30209 20085 30243
rect 20119 30209 20131 30243
rect 20340 30240 20352 30249
rect 20307 30212 20352 30240
rect 20073 30203 20131 30209
rect 20340 30203 20352 30212
rect 20346 30200 20352 30203
rect 20404 30200 20410 30252
rect 22554 30200 22560 30252
rect 22612 30240 22618 30252
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 22612 30212 23397 30240
rect 22612 30200 22618 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 19334 30172 19340 30184
rect 18892 30144 19340 30172
rect 19334 30132 19340 30144
rect 19392 30132 19398 30184
rect 23290 30172 23296 30184
rect 23251 30144 23296 30172
rect 23290 30132 23296 30144
rect 23348 30132 23354 30184
rect 24578 30132 24584 30184
rect 24636 30172 24642 30184
rect 24673 30175 24731 30181
rect 24673 30172 24685 30175
rect 24636 30144 24685 30172
rect 24636 30132 24642 30144
rect 24673 30141 24685 30144
rect 24719 30141 24731 30175
rect 25038 30172 25044 30184
rect 24999 30144 25044 30172
rect 24673 30135 24731 30141
rect 25038 30132 25044 30144
rect 25096 30132 25102 30184
rect 25133 30175 25191 30181
rect 25133 30141 25145 30175
rect 25179 30141 25191 30175
rect 25133 30135 25191 30141
rect 15838 30104 15844 30116
rect 14292 30076 15844 30104
rect 15838 30064 15844 30076
rect 15896 30064 15902 30116
rect 22278 30104 22284 30116
rect 22239 30076 22284 30104
rect 22278 30064 22284 30076
rect 22336 30064 22342 30116
rect 25148 30104 25176 30135
rect 25056 30076 25176 30104
rect 25056 30048 25084 30076
rect 10962 30036 10968 30048
rect 10428 30008 10968 30036
rect 9309 29999 9367 30005
rect 10962 29996 10968 30008
rect 11020 29996 11026 30048
rect 11057 30039 11115 30045
rect 11057 30005 11069 30039
rect 11103 30036 11115 30039
rect 12618 30036 12624 30048
rect 11103 30008 12624 30036
rect 11103 30005 11115 30008
rect 11057 29999 11115 30005
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 14458 29996 14464 30048
rect 14516 30036 14522 30048
rect 14737 30039 14795 30045
rect 14737 30036 14749 30039
rect 14516 30008 14749 30036
rect 14516 29996 14522 30008
rect 14737 30005 14749 30008
rect 14783 30005 14795 30039
rect 14737 29999 14795 30005
rect 15286 29996 15292 30048
rect 15344 30036 15350 30048
rect 15746 30036 15752 30048
rect 15344 30008 15752 30036
rect 15344 29996 15350 30008
rect 15746 29996 15752 30008
rect 15804 29996 15810 30048
rect 16117 30039 16175 30045
rect 16117 30005 16129 30039
rect 16163 30036 16175 30039
rect 16482 30036 16488 30048
rect 16163 30008 16488 30036
rect 16163 30005 16175 30008
rect 16117 29999 16175 30005
rect 16482 29996 16488 30008
rect 16540 29996 16546 30048
rect 17126 29996 17132 30048
rect 17184 30036 17190 30048
rect 18233 30039 18291 30045
rect 18233 30036 18245 30039
rect 17184 30008 18245 30036
rect 17184 29996 17190 30008
rect 18233 30005 18245 30008
rect 18279 30005 18291 30039
rect 21450 30036 21456 30048
rect 21411 30008 21456 30036
rect 18233 29999 18291 30005
rect 21450 29996 21456 30008
rect 21508 29996 21514 30048
rect 25038 29996 25044 30048
rect 25096 29996 25102 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 2593 29835 2651 29841
rect 2593 29801 2605 29835
rect 2639 29832 2651 29835
rect 2682 29832 2688 29844
rect 2639 29804 2688 29832
rect 2639 29801 2651 29804
rect 2593 29795 2651 29801
rect 2682 29792 2688 29804
rect 2740 29792 2746 29844
rect 3329 29835 3387 29841
rect 3329 29801 3341 29835
rect 3375 29832 3387 29835
rect 4062 29832 4068 29844
rect 3375 29804 4068 29832
rect 3375 29801 3387 29804
rect 3329 29795 3387 29801
rect 4062 29792 4068 29804
rect 4120 29792 4126 29844
rect 4154 29792 4160 29844
rect 4212 29832 4218 29844
rect 8018 29832 8024 29844
rect 4212 29804 8024 29832
rect 4212 29792 4218 29804
rect 8018 29792 8024 29804
rect 8076 29832 8082 29844
rect 11238 29832 11244 29844
rect 8076 29804 11244 29832
rect 8076 29792 8082 29804
rect 11238 29792 11244 29804
rect 11296 29832 11302 29844
rect 12066 29832 12072 29844
rect 11296 29804 12072 29832
rect 11296 29792 11302 29804
rect 12066 29792 12072 29804
rect 12124 29792 12130 29844
rect 14366 29832 14372 29844
rect 12452 29804 14372 29832
rect 3988 29736 5488 29764
rect 3878 29696 3884 29708
rect 2608 29668 3884 29696
rect 2608 29637 2636 29668
rect 3878 29656 3884 29668
rect 3936 29656 3942 29708
rect 2593 29631 2651 29637
rect 2593 29597 2605 29631
rect 2639 29597 2651 29631
rect 2593 29591 2651 29597
rect 2682 29588 2688 29640
rect 2740 29628 2746 29640
rect 2777 29631 2835 29637
rect 2777 29628 2789 29631
rect 2740 29600 2789 29628
rect 2740 29588 2746 29600
rect 2777 29597 2789 29600
rect 2823 29597 2835 29631
rect 2777 29591 2835 29597
rect 3237 29631 3295 29637
rect 3237 29597 3249 29631
rect 3283 29597 3295 29631
rect 3237 29591 3295 29597
rect 3421 29631 3479 29637
rect 3421 29597 3433 29631
rect 3467 29628 3479 29631
rect 3988 29628 4016 29736
rect 5460 29708 5488 29736
rect 9214 29724 9220 29776
rect 9272 29764 9278 29776
rect 12452 29764 12480 29804
rect 14366 29792 14372 29804
rect 14424 29792 14430 29844
rect 14553 29835 14611 29841
rect 14553 29801 14565 29835
rect 14599 29832 14611 29835
rect 14642 29832 14648 29844
rect 14599 29804 14648 29832
rect 14599 29801 14611 29804
rect 14553 29795 14611 29801
rect 14642 29792 14648 29804
rect 14700 29792 14706 29844
rect 15010 29792 15016 29844
rect 15068 29832 15074 29844
rect 15470 29832 15476 29844
rect 15068 29804 15476 29832
rect 15068 29792 15074 29804
rect 15470 29792 15476 29804
rect 15528 29792 15534 29844
rect 16022 29832 16028 29844
rect 15983 29804 16028 29832
rect 16022 29792 16028 29804
rect 16080 29792 16086 29844
rect 16482 29792 16488 29844
rect 16540 29832 16546 29844
rect 18233 29835 18291 29841
rect 18233 29832 18245 29835
rect 16540 29804 18245 29832
rect 16540 29792 16546 29804
rect 18233 29801 18245 29804
rect 18279 29801 18291 29835
rect 18414 29832 18420 29844
rect 18375 29804 18420 29832
rect 18233 29795 18291 29801
rect 9272 29736 12480 29764
rect 9272 29724 9278 29736
rect 12526 29724 12532 29776
rect 12584 29764 12590 29776
rect 14734 29764 14740 29776
rect 12584 29736 12629 29764
rect 13556 29736 14740 29764
rect 12584 29724 12590 29736
rect 4249 29699 4307 29705
rect 4249 29665 4261 29699
rect 4295 29696 4307 29699
rect 4614 29696 4620 29708
rect 4295 29668 4620 29696
rect 4295 29665 4307 29668
rect 4249 29659 4307 29665
rect 4614 29656 4620 29668
rect 4672 29656 4678 29708
rect 5442 29656 5448 29708
rect 5500 29696 5506 29708
rect 5721 29699 5779 29705
rect 5721 29696 5733 29699
rect 5500 29668 5733 29696
rect 5500 29656 5506 29668
rect 5721 29665 5733 29668
rect 5767 29665 5779 29699
rect 5721 29659 5779 29665
rect 5813 29699 5871 29705
rect 5813 29665 5825 29699
rect 5859 29696 5871 29699
rect 5902 29696 5908 29708
rect 5859 29668 5908 29696
rect 5859 29665 5871 29668
rect 5813 29659 5871 29665
rect 5902 29656 5908 29668
rect 5960 29656 5966 29708
rect 8110 29656 8116 29708
rect 8168 29696 8174 29708
rect 10318 29696 10324 29708
rect 8168 29668 10324 29696
rect 8168 29656 8174 29668
rect 10318 29656 10324 29668
rect 10376 29656 10382 29708
rect 10502 29656 10508 29708
rect 10560 29696 10566 29708
rect 12066 29696 12072 29708
rect 10560 29668 10732 29696
rect 12027 29668 12072 29696
rect 10560 29656 10566 29668
rect 3467 29600 4016 29628
rect 4157 29631 4215 29637
rect 3467 29597 3479 29600
rect 3421 29591 3479 29597
rect 4157 29597 4169 29631
rect 4203 29628 4215 29631
rect 5350 29628 5356 29640
rect 4203 29600 5356 29628
rect 4203 29597 4215 29600
rect 4157 29591 4215 29597
rect 3252 29492 3280 29591
rect 5350 29588 5356 29600
rect 5408 29588 5414 29640
rect 5534 29628 5540 29640
rect 5495 29600 5540 29628
rect 5534 29588 5540 29600
rect 5592 29588 5598 29640
rect 5629 29631 5687 29637
rect 5629 29597 5641 29631
rect 5675 29597 5687 29631
rect 5629 29591 5687 29597
rect 4798 29560 4804 29572
rect 4540 29532 4804 29560
rect 4540 29501 4568 29532
rect 4798 29520 4804 29532
rect 4856 29560 4862 29572
rect 5644 29560 5672 29591
rect 7282 29588 7288 29640
rect 7340 29628 7346 29640
rect 8202 29628 8208 29640
rect 7340 29600 8208 29628
rect 7340 29588 7346 29600
rect 8202 29588 8208 29600
rect 8260 29588 8266 29640
rect 9122 29628 9128 29640
rect 9083 29600 9128 29628
rect 9122 29588 9128 29600
rect 9180 29588 9186 29640
rect 9306 29588 9312 29640
rect 9364 29637 9370 29640
rect 9364 29631 9386 29637
rect 9374 29597 9386 29631
rect 9364 29591 9386 29597
rect 9493 29631 9551 29637
rect 9493 29597 9505 29631
rect 9539 29628 9551 29631
rect 9582 29628 9588 29640
rect 9539 29600 9588 29628
rect 9539 29597 9551 29600
rect 9493 29591 9551 29597
rect 9364 29588 9370 29591
rect 9582 29588 9588 29600
rect 9640 29588 9646 29640
rect 10704 29637 10732 29668
rect 12066 29656 12072 29668
rect 12124 29656 12130 29708
rect 13556 29696 13584 29736
rect 14734 29724 14740 29736
rect 14792 29764 14798 29776
rect 15286 29764 15292 29776
rect 14792 29736 15292 29764
rect 14792 29724 14798 29736
rect 15286 29724 15292 29736
rect 15344 29724 15350 29776
rect 18248 29764 18276 29795
rect 18414 29792 18420 29804
rect 18472 29792 18478 29844
rect 20349 29835 20407 29841
rect 20349 29801 20361 29835
rect 20395 29801 20407 29835
rect 20349 29795 20407 29801
rect 20364 29764 20392 29795
rect 20438 29792 20444 29844
rect 20496 29832 20502 29844
rect 20533 29835 20591 29841
rect 20533 29832 20545 29835
rect 20496 29804 20545 29832
rect 20496 29792 20502 29804
rect 20533 29801 20545 29804
rect 20579 29801 20591 29835
rect 21174 29832 21180 29844
rect 21135 29804 21180 29832
rect 20533 29795 20591 29801
rect 21174 29792 21180 29804
rect 21232 29792 21238 29844
rect 22741 29835 22799 29841
rect 22741 29801 22753 29835
rect 22787 29801 22799 29835
rect 22741 29795 22799 29801
rect 22925 29835 22983 29841
rect 22925 29801 22937 29835
rect 22971 29832 22983 29835
rect 23382 29832 23388 29844
rect 22971 29804 23388 29832
rect 22971 29801 22983 29804
rect 22925 29795 22983 29801
rect 18248 29736 20392 29764
rect 22756 29764 22784 29795
rect 23382 29792 23388 29804
rect 23440 29792 23446 29844
rect 24765 29835 24823 29841
rect 24765 29801 24777 29835
rect 24811 29832 24823 29835
rect 24854 29832 24860 29844
rect 24811 29804 24860 29832
rect 24811 29801 24823 29804
rect 24765 29795 24823 29801
rect 24854 29792 24860 29804
rect 24912 29792 24918 29844
rect 23290 29764 23296 29776
rect 22756 29736 23296 29764
rect 23290 29724 23296 29736
rect 23348 29724 23354 29776
rect 12176 29668 13584 29696
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29597 10655 29631
rect 10597 29591 10655 29597
rect 10689 29631 10747 29637
rect 10689 29597 10701 29631
rect 10735 29597 10747 29631
rect 10689 29591 10747 29597
rect 6822 29560 6828 29572
rect 4856 29532 5672 29560
rect 6380 29532 6828 29560
rect 4856 29520 4862 29532
rect 4525 29495 4583 29501
rect 4525 29492 4537 29495
rect 3252 29464 4537 29492
rect 4525 29461 4537 29464
rect 4571 29461 4583 29495
rect 4525 29455 4583 29461
rect 5353 29495 5411 29501
rect 5353 29461 5365 29495
rect 5399 29492 5411 29495
rect 6380 29492 6408 29532
rect 6822 29520 6828 29532
rect 6880 29520 6886 29572
rect 7006 29560 7012 29572
rect 6967 29532 7012 29560
rect 7006 29520 7012 29532
rect 7064 29520 7070 29572
rect 8389 29563 8447 29569
rect 8389 29529 8401 29563
rect 8435 29560 8447 29563
rect 8754 29560 8760 29572
rect 8435 29532 8760 29560
rect 8435 29529 8447 29532
rect 8389 29523 8447 29529
rect 8754 29520 8760 29532
rect 8812 29520 8818 29572
rect 10612 29560 10640 29591
rect 10778 29588 10784 29640
rect 10836 29628 10842 29640
rect 10836 29600 10881 29628
rect 10836 29588 10842 29600
rect 10962 29588 10968 29640
rect 11020 29628 11026 29640
rect 12176 29637 12204 29668
rect 13630 29656 13636 29708
rect 13688 29696 13694 29708
rect 17865 29699 17923 29705
rect 13688 29668 14412 29696
rect 13688 29656 13694 29668
rect 12161 29631 12219 29637
rect 11020 29600 12020 29628
rect 11020 29588 11026 29600
rect 11882 29560 11888 29572
rect 10612 29532 11888 29560
rect 11882 29520 11888 29532
rect 11940 29520 11946 29572
rect 7190 29492 7196 29504
rect 5399 29464 6408 29492
rect 7151 29464 7196 29492
rect 5399 29461 5411 29464
rect 5353 29455 5411 29461
rect 7190 29452 7196 29464
rect 7248 29452 7254 29504
rect 8570 29492 8576 29504
rect 8483 29464 8576 29492
rect 8570 29452 8576 29464
rect 8628 29492 8634 29504
rect 9217 29495 9275 29501
rect 9217 29492 9229 29495
rect 8628 29464 9229 29492
rect 8628 29452 8634 29464
rect 9217 29461 9229 29464
rect 9263 29461 9275 29495
rect 9217 29455 9275 29461
rect 9490 29452 9496 29504
rect 9548 29492 9554 29504
rect 10321 29495 10379 29501
rect 9548 29464 9593 29492
rect 9548 29452 9554 29464
rect 10321 29461 10333 29495
rect 10367 29492 10379 29495
rect 10686 29492 10692 29504
rect 10367 29464 10692 29492
rect 10367 29461 10379 29464
rect 10321 29455 10379 29461
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 11992 29492 12020 29600
rect 12161 29597 12173 29631
rect 12207 29597 12219 29631
rect 12161 29591 12219 29597
rect 12342 29588 12348 29640
rect 12400 29628 12406 29640
rect 13078 29628 13084 29640
rect 12400 29600 13084 29628
rect 12400 29588 12406 29600
rect 13078 29588 13084 29600
rect 13136 29588 13142 29640
rect 13357 29631 13415 29637
rect 13357 29597 13369 29631
rect 13403 29628 13415 29631
rect 13722 29628 13728 29640
rect 13403 29600 13728 29628
rect 13403 29597 13415 29600
rect 13357 29591 13415 29597
rect 13722 29588 13728 29600
rect 13780 29588 13786 29640
rect 14384 29637 14412 29668
rect 17865 29665 17877 29699
rect 17911 29696 17923 29699
rect 19334 29696 19340 29708
rect 17911 29668 19340 29696
rect 17911 29665 17923 29668
rect 17865 29659 17923 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 14277 29631 14335 29637
rect 14277 29597 14289 29631
rect 14323 29597 14335 29631
rect 14277 29591 14335 29597
rect 14369 29631 14427 29637
rect 14369 29597 14381 29631
rect 14415 29628 14427 29631
rect 14550 29628 14556 29640
rect 14415 29600 14556 29628
rect 14415 29597 14427 29600
rect 14369 29591 14427 29597
rect 14292 29560 14320 29591
rect 14550 29588 14556 29600
rect 14608 29588 14614 29640
rect 14645 29631 14703 29637
rect 14645 29597 14657 29631
rect 14691 29628 14703 29631
rect 14734 29628 14740 29640
rect 14691 29600 14740 29628
rect 14691 29597 14703 29600
rect 14645 29591 14703 29597
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 15286 29588 15292 29640
rect 15344 29628 15350 29640
rect 15344 29600 15389 29628
rect 15344 29588 15350 29600
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 16209 29631 16267 29637
rect 16209 29628 16221 29631
rect 15804 29600 16221 29628
rect 15804 29588 15810 29600
rect 16209 29597 16221 29600
rect 16255 29597 16267 29631
rect 16482 29628 16488 29640
rect 16443 29600 16488 29628
rect 16209 29591 16267 29597
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 19981 29631 20039 29637
rect 19981 29597 19993 29631
rect 20027 29628 20039 29631
rect 22465 29631 22523 29637
rect 20027 29600 21588 29628
rect 20027 29597 20039 29600
rect 19981 29591 20039 29597
rect 15654 29560 15660 29572
rect 14292 29532 15660 29560
rect 15654 29520 15660 29532
rect 15712 29560 15718 29572
rect 16500 29560 16528 29588
rect 15712 29532 16528 29560
rect 20993 29563 21051 29569
rect 15712 29520 15718 29532
rect 20993 29529 21005 29563
rect 21039 29560 21051 29563
rect 21450 29560 21456 29572
rect 21039 29532 21456 29560
rect 21039 29529 21051 29532
rect 20993 29523 21051 29529
rect 21450 29520 21456 29532
rect 21508 29520 21514 29572
rect 21560 29504 21588 29600
rect 22465 29597 22477 29631
rect 22511 29628 22523 29631
rect 23014 29628 23020 29640
rect 22511 29600 23020 29628
rect 22511 29597 22523 29600
rect 22465 29591 22523 29597
rect 23014 29588 23020 29600
rect 23072 29588 23078 29640
rect 25038 29628 25044 29640
rect 24999 29600 25044 29628
rect 25038 29588 25044 29600
rect 25096 29588 25102 29640
rect 24765 29563 24823 29569
rect 24765 29529 24777 29563
rect 24811 29560 24823 29563
rect 25130 29560 25136 29572
rect 24811 29532 25136 29560
rect 24811 29529 24823 29532
rect 24765 29523 24823 29529
rect 25130 29520 25136 29532
rect 25188 29520 25194 29572
rect 12526 29492 12532 29504
rect 11992 29464 12532 29492
rect 12526 29452 12532 29464
rect 12584 29492 12590 29504
rect 13541 29495 13599 29501
rect 13541 29492 13553 29495
rect 12584 29464 13553 29492
rect 12584 29452 12590 29464
rect 13541 29461 13553 29464
rect 13587 29461 13599 29495
rect 14458 29492 14464 29504
rect 14419 29464 14464 29492
rect 13541 29455 13599 29461
rect 14458 29452 14464 29464
rect 14516 29452 14522 29504
rect 14550 29452 14556 29504
rect 14608 29492 14614 29504
rect 16298 29492 16304 29504
rect 14608 29464 16304 29492
rect 14608 29452 14614 29464
rect 16298 29452 16304 29464
rect 16356 29492 16362 29504
rect 16393 29495 16451 29501
rect 16393 29492 16405 29495
rect 16356 29464 16405 29492
rect 16356 29452 16362 29464
rect 16393 29461 16405 29464
rect 16439 29461 16451 29495
rect 16393 29455 16451 29461
rect 17862 29452 17868 29504
rect 17920 29492 17926 29504
rect 18233 29495 18291 29501
rect 18233 29492 18245 29495
rect 17920 29464 18245 29492
rect 17920 29452 17926 29464
rect 18233 29461 18245 29464
rect 18279 29461 18291 29495
rect 18233 29455 18291 29461
rect 20070 29452 20076 29504
rect 20128 29492 20134 29504
rect 20349 29495 20407 29501
rect 20349 29492 20361 29495
rect 20128 29464 20361 29492
rect 20128 29452 20134 29464
rect 20349 29461 20361 29464
rect 20395 29461 20407 29495
rect 20349 29455 20407 29461
rect 20530 29452 20536 29504
rect 20588 29492 20594 29504
rect 21193 29495 21251 29501
rect 21193 29492 21205 29495
rect 20588 29464 21205 29492
rect 20588 29452 20594 29464
rect 21193 29461 21205 29464
rect 21239 29461 21251 29495
rect 21193 29455 21251 29461
rect 21361 29495 21419 29501
rect 21361 29461 21373 29495
rect 21407 29492 21419 29495
rect 21542 29492 21548 29504
rect 21407 29464 21548 29492
rect 21407 29461 21419 29464
rect 21361 29455 21419 29461
rect 21542 29452 21548 29464
rect 21600 29452 21606 29504
rect 24670 29452 24676 29504
rect 24728 29492 24734 29504
rect 24949 29495 25007 29501
rect 24949 29492 24961 29495
rect 24728 29464 24961 29492
rect 24728 29452 24734 29464
rect 24949 29461 24961 29464
rect 24995 29461 25007 29495
rect 24949 29455 25007 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 7006 29248 7012 29300
rect 7064 29288 7070 29300
rect 7101 29291 7159 29297
rect 7101 29288 7113 29291
rect 7064 29260 7113 29288
rect 7064 29248 7070 29260
rect 7101 29257 7113 29260
rect 7147 29257 7159 29291
rect 7101 29251 7159 29257
rect 8386 29248 8392 29300
rect 8444 29288 8450 29300
rect 9033 29291 9091 29297
rect 9033 29288 9045 29291
rect 8444 29260 9045 29288
rect 8444 29248 8450 29260
rect 9033 29257 9045 29260
rect 9079 29257 9091 29291
rect 9033 29251 9091 29257
rect 10778 29248 10784 29300
rect 10836 29288 10842 29300
rect 11793 29291 11851 29297
rect 11793 29288 11805 29291
rect 10836 29260 11805 29288
rect 10836 29248 10842 29260
rect 11793 29257 11805 29260
rect 11839 29257 11851 29291
rect 11793 29251 11851 29257
rect 12345 29291 12403 29297
rect 12345 29257 12357 29291
rect 12391 29288 12403 29291
rect 13262 29288 13268 29300
rect 12391 29260 13268 29288
rect 12391 29257 12403 29260
rect 12345 29251 12403 29257
rect 13262 29248 13268 29260
rect 13320 29248 13326 29300
rect 14277 29291 14335 29297
rect 14277 29257 14289 29291
rect 14323 29257 14335 29291
rect 14277 29251 14335 29257
rect 8205 29223 8263 29229
rect 8205 29189 8217 29223
rect 8251 29220 8263 29223
rect 8570 29220 8576 29232
rect 8251 29192 8576 29220
rect 8251 29189 8263 29192
rect 8205 29183 8263 29189
rect 8570 29180 8576 29192
rect 8628 29180 8634 29232
rect 9306 29220 9312 29232
rect 8680 29192 9312 29220
rect 3510 29112 3516 29164
rect 3568 29152 3574 29164
rect 3973 29155 4031 29161
rect 3973 29152 3985 29155
rect 3568 29124 3985 29152
rect 3568 29112 3574 29124
rect 3973 29121 3985 29124
rect 4019 29121 4031 29155
rect 6730 29152 6736 29164
rect 6691 29124 6736 29152
rect 3973 29115 4031 29121
rect 6730 29112 6736 29124
rect 6788 29112 6794 29164
rect 8021 29155 8079 29161
rect 8021 29121 8033 29155
rect 8067 29121 8079 29155
rect 8294 29152 8300 29164
rect 8255 29124 8300 29152
rect 8021 29115 8079 29121
rect 4709 29087 4767 29093
rect 4709 29053 4721 29087
rect 4755 29084 4767 29087
rect 4890 29084 4896 29096
rect 4755 29056 4896 29084
rect 4755 29053 4767 29056
rect 4709 29047 4767 29053
rect 4890 29044 4896 29056
rect 4948 29044 4954 29096
rect 4985 29087 5043 29093
rect 4985 29053 4997 29087
rect 5031 29084 5043 29087
rect 5350 29084 5356 29096
rect 5031 29056 5356 29084
rect 5031 29053 5043 29056
rect 4985 29047 5043 29053
rect 5350 29044 5356 29056
rect 5408 29044 5414 29096
rect 6825 29087 6883 29093
rect 6825 29053 6837 29087
rect 6871 29053 6883 29087
rect 8036 29084 8064 29115
rect 8294 29112 8300 29124
rect 8352 29112 8358 29164
rect 8386 29112 8392 29164
rect 8444 29152 8450 29164
rect 8680 29152 8708 29192
rect 9306 29180 9312 29192
rect 9364 29180 9370 29232
rect 9490 29180 9496 29232
rect 9548 29180 9554 29232
rect 12618 29220 12624 29232
rect 12579 29192 12624 29220
rect 12618 29180 12624 29192
rect 12676 29180 12682 29232
rect 13538 29180 13544 29232
rect 13596 29220 13602 29232
rect 13725 29223 13783 29229
rect 13725 29220 13737 29223
rect 13596 29192 13737 29220
rect 13596 29180 13602 29192
rect 13725 29189 13737 29192
rect 13771 29189 13783 29223
rect 14292 29220 14320 29251
rect 15286 29248 15292 29300
rect 15344 29288 15350 29300
rect 16206 29288 16212 29300
rect 15344 29260 16212 29288
rect 15344 29248 15350 29260
rect 16206 29248 16212 29260
rect 16264 29288 16270 29300
rect 16301 29291 16359 29297
rect 16301 29288 16313 29291
rect 16264 29260 16313 29288
rect 16264 29248 16270 29260
rect 16301 29257 16313 29260
rect 16347 29257 16359 29291
rect 17862 29288 17868 29300
rect 17823 29260 17868 29288
rect 16301 29251 16359 29257
rect 17862 29248 17868 29260
rect 17920 29248 17926 29300
rect 20070 29288 20076 29300
rect 18800 29260 19104 29288
rect 20031 29260 20076 29288
rect 15166 29223 15224 29229
rect 15166 29220 15178 29223
rect 14292 29192 15178 29220
rect 13725 29183 13783 29189
rect 15166 29189 15178 29192
rect 15212 29189 15224 29223
rect 15166 29183 15224 29189
rect 15746 29180 15752 29232
rect 15804 29220 15810 29232
rect 17405 29223 17463 29229
rect 17405 29220 17417 29223
rect 15804 29192 17417 29220
rect 15804 29180 15810 29192
rect 17405 29189 17417 29192
rect 17451 29220 17463 29223
rect 17586 29220 17592 29232
rect 17451 29192 17592 29220
rect 17451 29189 17463 29192
rect 17405 29183 17463 29189
rect 17586 29180 17592 29192
rect 17644 29180 17650 29232
rect 18800 29229 18828 29260
rect 18785 29223 18843 29229
rect 18785 29220 18797 29223
rect 18064 29192 18797 29220
rect 8444 29124 8708 29152
rect 9217 29155 9275 29161
rect 8444 29112 8450 29124
rect 9217 29121 9229 29155
rect 9263 29152 9275 29155
rect 9508 29152 9536 29180
rect 10318 29152 10324 29164
rect 9263 29124 9536 29152
rect 10279 29124 10324 29152
rect 9263 29121 9275 29124
rect 9217 29115 9275 29121
rect 10318 29112 10324 29124
rect 10376 29112 10382 29164
rect 11698 29152 11704 29164
rect 11659 29124 11704 29152
rect 11698 29112 11704 29124
rect 11756 29112 11762 29164
rect 11882 29152 11888 29164
rect 11843 29124 11888 29152
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 12345 29155 12403 29161
rect 12345 29121 12357 29155
rect 12391 29152 12403 29155
rect 12434 29152 12440 29164
rect 12391 29124 12440 29152
rect 12391 29121 12403 29124
rect 12345 29115 12403 29121
rect 12434 29112 12440 29124
rect 12492 29112 12498 29164
rect 13633 29155 13691 29161
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13633 29115 13691 29121
rect 14461 29155 14519 29161
rect 14461 29121 14473 29155
rect 14507 29152 14519 29155
rect 14734 29152 14740 29164
rect 14507 29124 14740 29152
rect 14507 29121 14519 29124
rect 14461 29115 14519 29121
rect 8662 29084 8668 29096
rect 8036 29056 8668 29084
rect 6825 29047 6883 29053
rect 4154 29016 4160 29028
rect 4115 28988 4160 29016
rect 4154 28976 4160 28988
rect 4212 28976 4218 29028
rect 6840 29016 6868 29047
rect 8662 29044 8668 29056
rect 8720 29084 8726 29096
rect 9122 29084 9128 29096
rect 8720 29056 9128 29084
rect 8720 29044 8726 29056
rect 9122 29044 9128 29056
rect 9180 29044 9186 29096
rect 9309 29087 9367 29093
rect 9309 29053 9321 29087
rect 9355 29053 9367 29087
rect 9309 29047 9367 29053
rect 9401 29087 9459 29093
rect 9401 29053 9413 29087
rect 9447 29053 9459 29087
rect 9401 29047 9459 29053
rect 8478 29016 8484 29028
rect 6840 28988 8484 29016
rect 8478 28976 8484 28988
rect 8536 28976 8542 29028
rect 8573 29019 8631 29025
rect 8573 28985 8585 29019
rect 8619 29016 8631 29019
rect 9324 29016 9352 29047
rect 8619 28988 9352 29016
rect 9416 29016 9444 29047
rect 9490 29044 9496 29096
rect 9548 29084 9554 29096
rect 10594 29084 10600 29096
rect 9548 29056 9593 29084
rect 10555 29056 10600 29084
rect 9548 29044 9554 29056
rect 10594 29044 10600 29056
rect 10652 29044 10658 29096
rect 13648 29084 13676 29115
rect 14734 29112 14740 29124
rect 14792 29112 14798 29164
rect 14918 29152 14924 29164
rect 14879 29124 14924 29152
rect 14918 29112 14924 29124
rect 14976 29112 14982 29164
rect 16758 29152 16764 29164
rect 15028 29124 16764 29152
rect 15028 29084 15056 29124
rect 16758 29112 16764 29124
rect 16816 29112 16822 29164
rect 17126 29112 17132 29164
rect 17184 29152 17190 29164
rect 18064 29161 18092 29192
rect 18785 29189 18797 29192
rect 18831 29189 18843 29223
rect 18985 29223 19043 29229
rect 18985 29220 18997 29223
rect 18785 29183 18843 29189
rect 18892 29192 18997 29220
rect 17221 29155 17279 29161
rect 17221 29152 17233 29155
rect 17184 29124 17233 29152
rect 17184 29112 17190 29124
rect 17221 29121 17233 29124
rect 17267 29121 17279 29155
rect 17221 29115 17279 29121
rect 18049 29155 18107 29161
rect 18049 29121 18061 29155
rect 18095 29121 18107 29155
rect 18230 29152 18236 29164
rect 18191 29124 18236 29152
rect 18049 29115 18107 29121
rect 18230 29112 18236 29124
rect 18288 29112 18294 29164
rect 18325 29155 18383 29161
rect 18325 29121 18337 29155
rect 18371 29152 18383 29155
rect 18892 29152 18920 29192
rect 18985 29189 18997 29192
rect 19031 29189 19043 29223
rect 18985 29183 19043 29189
rect 18371 29124 18920 29152
rect 18371 29121 18383 29124
rect 18325 29115 18383 29121
rect 13648 29056 15056 29084
rect 17954 29044 17960 29096
rect 18012 29084 18018 29096
rect 18340 29084 18368 29115
rect 18012 29056 18368 29084
rect 19076 29084 19104 29260
rect 20070 29248 20076 29260
rect 20128 29248 20134 29300
rect 24857 29291 24915 29297
rect 24857 29257 24869 29291
rect 24903 29288 24915 29291
rect 25038 29288 25044 29300
rect 24903 29260 25044 29288
rect 24903 29257 24915 29260
rect 24857 29251 24915 29257
rect 25038 29248 25044 29260
rect 25096 29248 25102 29300
rect 19150 29180 19156 29232
rect 19208 29220 19214 29232
rect 20441 29223 20499 29229
rect 20441 29220 20453 29223
rect 19208 29192 20453 29220
rect 19208 29180 19214 29192
rect 20441 29189 20453 29192
rect 20487 29189 20499 29223
rect 20441 29183 20499 29189
rect 22005 29223 22063 29229
rect 22005 29189 22017 29223
rect 22051 29220 22063 29223
rect 22738 29220 22744 29232
rect 22051 29192 22744 29220
rect 22051 29189 22063 29192
rect 22005 29183 22063 29189
rect 22738 29180 22744 29192
rect 22796 29180 22802 29232
rect 20257 29155 20315 29161
rect 20257 29121 20269 29155
rect 20303 29121 20315 29155
rect 20530 29152 20536 29164
rect 20491 29124 20536 29152
rect 20257 29115 20315 29121
rect 19426 29084 19432 29096
rect 19076 29056 19432 29084
rect 18012 29044 18018 29056
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 20272 29084 20300 29115
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 20898 29112 20904 29164
rect 20956 29152 20962 29164
rect 20993 29155 21051 29161
rect 20993 29152 21005 29155
rect 20956 29124 21005 29152
rect 20956 29112 20962 29124
rect 20993 29121 21005 29124
rect 21039 29121 21051 29155
rect 21174 29152 21180 29164
rect 21135 29124 21180 29152
rect 20993 29115 21051 29121
rect 21174 29112 21180 29124
rect 21232 29112 21238 29164
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29152 21327 29155
rect 21450 29152 21456 29164
rect 21315 29124 21456 29152
rect 21315 29121 21327 29124
rect 21269 29115 21327 29121
rect 21284 29084 21312 29115
rect 21450 29112 21456 29124
rect 21508 29112 21514 29164
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 22152 29124 22201 29152
rect 22152 29112 22158 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 23017 29155 23075 29161
rect 23017 29121 23029 29155
rect 23063 29152 23075 29155
rect 23106 29152 23112 29164
rect 23063 29124 23112 29152
rect 23063 29121 23075 29124
rect 23017 29115 23075 29121
rect 23106 29112 23112 29124
rect 23164 29112 23170 29164
rect 24489 29155 24547 29161
rect 24489 29152 24501 29155
rect 23400 29124 24501 29152
rect 22922 29084 22928 29096
rect 20272 29056 21312 29084
rect 22883 29056 22928 29084
rect 22922 29044 22928 29056
rect 22980 29044 22986 29096
rect 10962 29016 10968 29028
rect 9416 28988 10968 29016
rect 8619 28985 8631 28988
rect 8573 28979 8631 28985
rect 10962 28976 10968 28988
rect 11020 28976 11026 29028
rect 12250 28976 12256 29028
rect 12308 29016 12314 29028
rect 12437 29019 12495 29025
rect 12437 29016 12449 29019
rect 12308 28988 12449 29016
rect 12308 28976 12314 28988
rect 12437 28985 12449 28988
rect 12483 28985 12495 29019
rect 19153 29019 19211 29025
rect 12437 28979 12495 28985
rect 13648 28988 13860 29016
rect 8294 28908 8300 28960
rect 8352 28948 8358 28960
rect 9582 28948 9588 28960
rect 8352 28920 9588 28948
rect 8352 28908 8358 28920
rect 9582 28908 9588 28920
rect 9640 28908 9646 28960
rect 11882 28908 11888 28960
rect 11940 28948 11946 28960
rect 13648 28948 13676 28988
rect 11940 28920 13676 28948
rect 13832 28948 13860 28988
rect 16224 28988 16436 29016
rect 16224 28948 16252 28988
rect 13832 28920 16252 28948
rect 16408 28948 16436 28988
rect 17236 28988 17448 29016
rect 17236 28948 17264 28988
rect 16408 28920 17264 28948
rect 17420 28948 17448 28988
rect 19153 28985 19165 29019
rect 19199 29016 19211 29019
rect 19334 29016 19340 29028
rect 19199 28988 19340 29016
rect 19199 28985 19211 28988
rect 19153 28979 19211 28985
rect 19334 28976 19340 28988
rect 19392 29016 19398 29028
rect 20530 29016 20536 29028
rect 19392 28988 20536 29016
rect 19392 28976 19398 28988
rect 20530 28976 20536 28988
rect 20588 28976 20594 29028
rect 23400 29025 23428 29124
rect 24489 29121 24501 29124
rect 24535 29121 24547 29155
rect 24489 29115 24547 29121
rect 24581 29087 24639 29093
rect 24581 29053 24593 29087
rect 24627 29084 24639 29087
rect 25038 29084 25044 29096
rect 24627 29056 25044 29084
rect 24627 29053 24639 29056
rect 24581 29047 24639 29053
rect 25038 29044 25044 29056
rect 25096 29044 25102 29096
rect 23385 29019 23443 29025
rect 23385 28985 23397 29019
rect 23431 28985 23443 29019
rect 23385 28979 23443 28985
rect 18230 28948 18236 28960
rect 17420 28920 18236 28948
rect 11940 28908 11946 28920
rect 18230 28908 18236 28920
rect 18288 28948 18294 28960
rect 18969 28951 19027 28957
rect 18969 28948 18981 28951
rect 18288 28920 18981 28948
rect 18288 28908 18294 28920
rect 18969 28917 18981 28920
rect 19015 28917 19027 28951
rect 20990 28948 20996 28960
rect 20951 28920 20996 28948
rect 18969 28911 19027 28917
rect 20990 28908 20996 28920
rect 21048 28908 21054 28960
rect 22370 28948 22376 28960
rect 22331 28920 22376 28948
rect 22370 28908 22376 28920
rect 22428 28908 22434 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 4433 28747 4491 28753
rect 4433 28713 4445 28747
rect 4479 28744 4491 28747
rect 4890 28744 4896 28756
rect 4479 28716 4896 28744
rect 4479 28713 4491 28716
rect 4433 28707 4491 28713
rect 4890 28704 4896 28716
rect 4948 28744 4954 28756
rect 4948 28716 5212 28744
rect 4948 28704 4954 28716
rect 4154 28540 4160 28552
rect 4115 28512 4160 28540
rect 4154 28500 4160 28512
rect 4212 28500 4218 28552
rect 5184 28549 5212 28716
rect 5258 28704 5264 28756
rect 5316 28744 5322 28756
rect 5445 28747 5503 28753
rect 5445 28744 5457 28747
rect 5316 28716 5457 28744
rect 5316 28704 5322 28716
rect 5445 28713 5457 28716
rect 5491 28744 5503 28747
rect 5491 28716 6316 28744
rect 5491 28713 5503 28716
rect 5445 28707 5503 28713
rect 5169 28543 5227 28549
rect 5169 28509 5181 28543
rect 5215 28540 5227 28543
rect 5350 28540 5356 28552
rect 5215 28512 5356 28540
rect 5215 28509 5227 28512
rect 5169 28503 5227 28509
rect 5350 28500 5356 28512
rect 5408 28540 5414 28552
rect 6181 28543 6239 28549
rect 6181 28540 6193 28543
rect 5408 28512 6193 28540
rect 5408 28500 5414 28512
rect 6181 28509 6193 28512
rect 6227 28509 6239 28543
rect 6181 28503 6239 28509
rect 3970 28364 3976 28416
rect 4028 28404 4034 28416
rect 4617 28407 4675 28413
rect 4617 28404 4629 28407
rect 4028 28376 4629 28404
rect 4028 28364 4034 28376
rect 4617 28373 4629 28376
rect 4663 28373 4675 28407
rect 4617 28367 4675 28373
rect 5258 28364 5264 28416
rect 5316 28404 5322 28416
rect 5629 28407 5687 28413
rect 5629 28404 5641 28407
rect 5316 28376 5641 28404
rect 5316 28364 5322 28376
rect 5629 28373 5641 28376
rect 5675 28373 5687 28407
rect 6288 28404 6316 28716
rect 7466 28704 7472 28756
rect 7524 28744 7530 28756
rect 7561 28747 7619 28753
rect 7561 28744 7573 28747
rect 7524 28716 7573 28744
rect 7524 28704 7530 28716
rect 7561 28713 7573 28716
rect 7607 28713 7619 28747
rect 8386 28744 8392 28756
rect 7561 28707 7619 28713
rect 7852 28716 8392 28744
rect 6914 28636 6920 28688
rect 6972 28636 6978 28688
rect 7009 28679 7067 28685
rect 7009 28645 7021 28679
rect 7055 28676 7067 28679
rect 7852 28676 7880 28716
rect 8386 28704 8392 28716
rect 8444 28704 8450 28756
rect 8754 28704 8760 28756
rect 8812 28744 8818 28756
rect 9398 28744 9404 28756
rect 8812 28716 9404 28744
rect 8812 28704 8818 28716
rect 9398 28704 9404 28716
rect 9456 28704 9462 28756
rect 9582 28744 9588 28756
rect 9543 28716 9588 28744
rect 9582 28704 9588 28716
rect 9640 28704 9646 28756
rect 11882 28704 11888 28756
rect 11940 28744 11946 28756
rect 11977 28747 12035 28753
rect 11977 28744 11989 28747
rect 11940 28716 11989 28744
rect 11940 28704 11946 28716
rect 11977 28713 11989 28716
rect 12023 28713 12035 28747
rect 11977 28707 12035 28713
rect 14274 28704 14280 28756
rect 14332 28744 14338 28756
rect 15473 28747 15531 28753
rect 15473 28744 15485 28747
rect 14332 28716 15485 28744
rect 14332 28704 14338 28716
rect 15473 28713 15485 28716
rect 15519 28744 15531 28747
rect 16209 28747 16267 28753
rect 16209 28744 16221 28747
rect 15519 28716 16221 28744
rect 15519 28713 15531 28716
rect 15473 28707 15531 28713
rect 16209 28713 16221 28716
rect 16255 28744 16267 28747
rect 17034 28744 17040 28756
rect 16255 28716 17040 28744
rect 16255 28713 16267 28716
rect 16209 28707 16267 28713
rect 17034 28704 17040 28716
rect 17092 28704 17098 28756
rect 25038 28744 25044 28756
rect 24999 28716 25044 28744
rect 25038 28704 25044 28716
rect 25096 28704 25102 28756
rect 7055 28648 7880 28676
rect 7055 28645 7067 28648
rect 7009 28639 7067 28645
rect 6932 28608 6960 28636
rect 6932 28580 7052 28608
rect 6822 28500 6828 28552
rect 6880 28540 6886 28552
rect 6917 28543 6975 28549
rect 6917 28540 6929 28543
rect 6880 28512 6929 28540
rect 6880 28500 6886 28512
rect 6917 28509 6929 28512
rect 6963 28509 6975 28543
rect 7024 28540 7052 28580
rect 7190 28568 7196 28620
rect 7248 28608 7254 28620
rect 7852 28617 7880 28648
rect 14642 28636 14648 28688
rect 14700 28636 14706 28688
rect 15381 28679 15439 28685
rect 15381 28645 15393 28679
rect 15427 28676 15439 28679
rect 18322 28676 18328 28688
rect 15427 28648 18328 28676
rect 15427 28645 15439 28648
rect 15381 28639 15439 28645
rect 18322 28636 18328 28648
rect 18380 28636 18386 28688
rect 18782 28676 18788 28688
rect 18743 28648 18788 28676
rect 18782 28636 18788 28648
rect 18840 28676 18846 28688
rect 19058 28676 19064 28688
rect 18840 28648 19064 28676
rect 18840 28636 18846 28648
rect 19058 28636 19064 28648
rect 19116 28636 19122 28688
rect 19429 28679 19487 28685
rect 19429 28645 19441 28679
rect 19475 28676 19487 28679
rect 20898 28676 20904 28688
rect 19475 28648 20904 28676
rect 19475 28645 19487 28648
rect 19429 28639 19487 28645
rect 20898 28636 20904 28648
rect 20956 28676 20962 28688
rect 21453 28679 21511 28685
rect 20956 28648 21128 28676
rect 20956 28636 20962 28648
rect 7745 28611 7803 28617
rect 7745 28608 7757 28611
rect 7248 28580 7757 28608
rect 7248 28568 7254 28580
rect 7745 28577 7757 28580
rect 7791 28577 7803 28611
rect 7745 28571 7803 28577
rect 7837 28611 7895 28617
rect 7837 28577 7849 28611
rect 7883 28577 7895 28611
rect 10502 28608 10508 28620
rect 7837 28571 7895 28577
rect 7944 28580 10508 28608
rect 7101 28543 7159 28549
rect 7101 28540 7113 28543
rect 7024 28512 7113 28540
rect 6917 28503 6975 28509
rect 7101 28509 7113 28512
rect 7147 28509 7159 28543
rect 7101 28503 7159 28509
rect 7282 28500 7288 28552
rect 7340 28540 7346 28552
rect 7944 28549 7972 28580
rect 10502 28568 10508 28580
rect 10560 28568 10566 28620
rect 14660 28608 14688 28636
rect 14292 28580 14688 28608
rect 7929 28543 7987 28549
rect 7929 28540 7941 28543
rect 7340 28512 7941 28540
rect 7340 28500 7346 28512
rect 7929 28509 7941 28512
rect 7975 28509 7987 28543
rect 7929 28503 7987 28509
rect 8018 28500 8024 28552
rect 8076 28540 8082 28552
rect 8076 28512 8121 28540
rect 8076 28500 8082 28512
rect 8478 28500 8484 28552
rect 8536 28540 8542 28552
rect 9125 28543 9183 28549
rect 9125 28540 9137 28543
rect 8536 28512 9137 28540
rect 8536 28500 8542 28512
rect 9125 28509 9137 28512
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 9674 28500 9680 28552
rect 9732 28540 9738 28552
rect 10594 28540 10600 28552
rect 9732 28512 10600 28540
rect 9732 28500 9738 28512
rect 10594 28500 10600 28512
rect 10652 28500 10658 28552
rect 10686 28500 10692 28552
rect 10744 28540 10750 28552
rect 14292 28549 14320 28580
rect 14734 28568 14740 28620
rect 14792 28608 14798 28620
rect 16574 28608 16580 28620
rect 14792 28580 14837 28608
rect 16040 28580 16580 28608
rect 14792 28568 14798 28580
rect 10853 28543 10911 28549
rect 10853 28540 10865 28543
rect 10744 28512 10865 28540
rect 10744 28500 10750 28512
rect 10853 28509 10865 28512
rect 10899 28509 10911 28543
rect 10853 28503 10911 28509
rect 14277 28543 14335 28549
rect 14277 28509 14289 28543
rect 14323 28509 14335 28543
rect 14550 28540 14556 28552
rect 14511 28512 14556 28540
rect 14277 28503 14335 28509
rect 14550 28500 14556 28512
rect 14608 28500 14614 28552
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28509 14703 28543
rect 14645 28503 14703 28509
rect 6365 28475 6423 28481
rect 6365 28441 6377 28475
rect 6411 28472 6423 28475
rect 6730 28472 6736 28484
rect 6411 28444 6736 28472
rect 6411 28441 6423 28444
rect 6365 28435 6423 28441
rect 6730 28432 6736 28444
rect 6788 28472 6794 28484
rect 8754 28472 8760 28484
rect 6788 28444 8760 28472
rect 6788 28432 6794 28444
rect 8754 28432 8760 28444
rect 8812 28432 8818 28484
rect 12802 28432 12808 28484
rect 12860 28472 12866 28484
rect 14660 28472 14688 28503
rect 15010 28500 15016 28552
rect 15068 28540 15074 28552
rect 15378 28540 15384 28552
rect 15068 28512 15384 28540
rect 15068 28500 15074 28512
rect 15378 28500 15384 28512
rect 15436 28540 15442 28552
rect 16040 28549 16068 28580
rect 16574 28568 16580 28580
rect 16632 28608 16638 28620
rect 16758 28608 16764 28620
rect 16632 28580 16764 28608
rect 16632 28568 16638 28580
rect 16758 28568 16764 28580
rect 16816 28568 16822 28620
rect 18877 28611 18935 28617
rect 18877 28577 18889 28611
rect 18923 28608 18935 28611
rect 19889 28611 19947 28617
rect 19889 28608 19901 28611
rect 18923 28580 19901 28608
rect 18923 28577 18935 28580
rect 18877 28571 18935 28577
rect 19889 28577 19901 28580
rect 19935 28577 19947 28611
rect 19889 28571 19947 28577
rect 20714 28568 20720 28620
rect 20772 28608 20778 28620
rect 20993 28611 21051 28617
rect 20993 28608 21005 28611
rect 20772 28580 21005 28608
rect 20772 28568 20778 28580
rect 20993 28577 21005 28580
rect 21039 28577 21051 28611
rect 20993 28571 21051 28577
rect 15565 28543 15623 28549
rect 15565 28540 15577 28543
rect 15436 28512 15577 28540
rect 15436 28500 15442 28512
rect 15565 28509 15577 28512
rect 15611 28509 15623 28543
rect 15565 28503 15623 28509
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 16117 28543 16175 28549
rect 16117 28509 16129 28543
rect 16163 28509 16175 28543
rect 16117 28503 16175 28509
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28540 17831 28543
rect 17954 28540 17960 28552
rect 17819 28512 17960 28540
rect 17819 28509 17831 28512
rect 17773 28503 17831 28509
rect 15194 28472 15200 28484
rect 12860 28444 14688 28472
rect 15155 28444 15200 28472
rect 12860 28432 12866 28444
rect 15194 28432 15200 28444
rect 15252 28432 15258 28484
rect 15580 28472 15608 28503
rect 16132 28472 16160 28503
rect 17954 28500 17960 28512
rect 18012 28500 18018 28552
rect 18966 28500 18972 28552
rect 19024 28540 19030 28552
rect 21100 28549 21128 28648
rect 21453 28645 21465 28679
rect 21499 28676 21511 28679
rect 22922 28676 22928 28688
rect 21499 28648 22928 28676
rect 21499 28645 21511 28648
rect 21453 28639 21511 28645
rect 22922 28636 22928 28648
rect 22980 28636 22986 28688
rect 23477 28679 23535 28685
rect 23477 28645 23489 28679
rect 23523 28676 23535 28679
rect 23523 28648 24716 28676
rect 23523 28645 23535 28648
rect 23477 28639 23535 28645
rect 23014 28608 23020 28620
rect 22975 28580 23020 28608
rect 23014 28568 23020 28580
rect 23072 28568 23078 28620
rect 24688 28617 24716 28648
rect 24673 28611 24731 28617
rect 24673 28577 24685 28611
rect 24719 28577 24731 28611
rect 24673 28571 24731 28577
rect 19613 28543 19671 28549
rect 19613 28540 19625 28543
rect 19024 28512 19625 28540
rect 19024 28500 19030 28512
rect 19613 28509 19625 28512
rect 19659 28509 19671 28543
rect 19613 28503 19671 28509
rect 19705 28543 19763 28549
rect 19705 28509 19717 28543
rect 19751 28509 19763 28543
rect 19705 28503 19763 28509
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28509 21143 28543
rect 22186 28540 22192 28552
rect 22147 28512 22192 28540
rect 21085 28503 21143 28509
rect 15580 28444 16160 28472
rect 18138 28432 18144 28484
rect 18196 28472 18202 28484
rect 18417 28475 18475 28481
rect 18417 28472 18429 28475
rect 18196 28444 18429 28472
rect 18196 28432 18202 28444
rect 18417 28441 18429 28444
rect 18463 28441 18475 28475
rect 18417 28435 18475 28441
rect 19426 28432 19432 28484
rect 19484 28472 19490 28484
rect 19720 28472 19748 28503
rect 19484 28444 19748 28472
rect 19484 28432 19490 28444
rect 11790 28404 11796 28416
rect 6288 28376 11796 28404
rect 5629 28367 5687 28373
rect 11790 28364 11796 28376
rect 11848 28364 11854 28416
rect 14369 28407 14427 28413
rect 14369 28373 14381 28407
rect 14415 28404 14427 28407
rect 14642 28404 14648 28416
rect 14415 28376 14648 28404
rect 14415 28373 14427 28376
rect 14369 28367 14427 28373
rect 14642 28364 14648 28376
rect 14700 28364 14706 28416
rect 15286 28404 15292 28416
rect 15247 28376 15292 28404
rect 15286 28364 15292 28376
rect 15344 28364 15350 28416
rect 16390 28404 16396 28416
rect 16351 28376 16396 28404
rect 16390 28364 16396 28376
rect 16448 28364 16454 28416
rect 17218 28364 17224 28416
rect 17276 28404 17282 28416
rect 17865 28407 17923 28413
rect 17865 28404 17877 28407
rect 17276 28376 17877 28404
rect 17276 28364 17282 28376
rect 17865 28373 17877 28376
rect 17911 28404 17923 28407
rect 19812 28404 19840 28503
rect 22186 28500 22192 28512
rect 22244 28500 22250 28552
rect 22370 28540 22376 28552
rect 22331 28512 22376 28540
rect 22370 28500 22376 28512
rect 22428 28500 22434 28552
rect 22465 28543 22523 28549
rect 22465 28509 22477 28543
rect 22511 28540 22523 28543
rect 23109 28543 23167 28549
rect 23109 28540 23121 28543
rect 22511 28512 23121 28540
rect 22511 28509 22523 28512
rect 22465 28503 22523 28509
rect 23109 28509 23121 28512
rect 23155 28540 23167 28543
rect 23198 28540 23204 28552
rect 23155 28512 23204 28540
rect 23155 28509 23167 28512
rect 23109 28503 23167 28509
rect 23198 28500 23204 28512
rect 23256 28500 23262 28552
rect 24302 28500 24308 28552
rect 24360 28540 24366 28552
rect 24765 28543 24823 28549
rect 24765 28540 24777 28543
rect 24360 28512 24777 28540
rect 24360 28500 24366 28512
rect 24765 28509 24777 28512
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 17911 28376 19840 28404
rect 22005 28407 22063 28413
rect 17911 28373 17923 28376
rect 17865 28367 17923 28373
rect 22005 28373 22017 28407
rect 22051 28404 22063 28407
rect 23106 28404 23112 28416
rect 22051 28376 23112 28404
rect 22051 28373 22063 28376
rect 22005 28367 22063 28373
rect 23106 28364 23112 28376
rect 23164 28364 23170 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 3510 28200 3516 28212
rect 3471 28172 3516 28200
rect 3510 28160 3516 28172
rect 3568 28200 3574 28212
rect 4614 28200 4620 28212
rect 3568 28172 4620 28200
rect 3568 28160 3574 28172
rect 4614 28160 4620 28172
rect 4672 28160 4678 28212
rect 5077 28203 5135 28209
rect 5077 28169 5089 28203
rect 5123 28200 5135 28203
rect 5350 28200 5356 28212
rect 5123 28172 5356 28200
rect 5123 28169 5135 28172
rect 5077 28163 5135 28169
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 5534 28160 5540 28212
rect 5592 28200 5598 28212
rect 5813 28203 5871 28209
rect 5813 28200 5825 28203
rect 5592 28172 5825 28200
rect 5592 28160 5598 28172
rect 5813 28169 5825 28172
rect 5859 28169 5871 28203
rect 5813 28163 5871 28169
rect 7834 28160 7840 28212
rect 7892 28209 7898 28212
rect 7892 28203 7911 28209
rect 7899 28169 7911 28203
rect 8018 28200 8024 28212
rect 7979 28172 8024 28200
rect 7892 28163 7911 28169
rect 7892 28160 7898 28163
rect 8018 28160 8024 28172
rect 8076 28160 8082 28212
rect 8662 28200 8668 28212
rect 8623 28172 8668 28200
rect 8662 28160 8668 28172
rect 8720 28160 8726 28212
rect 9490 28200 9496 28212
rect 9451 28172 9496 28200
rect 9490 28160 9496 28172
rect 9548 28160 9554 28212
rect 18690 28200 18696 28212
rect 12406 28172 18696 28200
rect 1670 28092 1676 28144
rect 1728 28132 1734 28144
rect 6086 28132 6092 28144
rect 1728 28104 6092 28132
rect 1728 28092 1734 28104
rect 6086 28092 6092 28104
rect 6144 28092 6150 28144
rect 7650 28132 7656 28144
rect 7611 28104 7656 28132
rect 7650 28092 7656 28104
rect 7708 28092 7714 28144
rect 9125 28135 9183 28141
rect 9125 28132 9137 28135
rect 8220 28104 9137 28132
rect 2406 28073 2412 28076
rect 2400 28027 2412 28073
rect 2464 28064 2470 28076
rect 3970 28064 3976 28076
rect 2464 28036 2500 28064
rect 3931 28036 3976 28064
rect 2406 28024 2412 28027
rect 2464 28024 2470 28036
rect 3970 28024 3976 28036
rect 4028 28024 4034 28076
rect 4157 28067 4215 28073
rect 4157 28033 4169 28067
rect 4203 28064 4215 28067
rect 5261 28067 5319 28073
rect 5261 28064 5273 28067
rect 4203 28036 5273 28064
rect 4203 28033 4215 28036
rect 4157 28027 4215 28033
rect 5261 28033 5273 28036
rect 5307 28064 5319 28067
rect 5626 28064 5632 28076
rect 5307 28036 5632 28064
rect 5307 28033 5319 28036
rect 5261 28027 5319 28033
rect 5626 28024 5632 28036
rect 5684 28024 5690 28076
rect 5718 28024 5724 28076
rect 5776 28064 5782 28076
rect 7668 28064 7696 28092
rect 8220 28064 8248 28104
rect 9125 28101 9137 28104
rect 9171 28101 9183 28135
rect 9125 28095 9183 28101
rect 9341 28135 9399 28141
rect 9341 28101 9353 28135
rect 9387 28132 9399 28135
rect 9858 28132 9864 28144
rect 9387 28104 9864 28132
rect 9387 28101 9399 28104
rect 9341 28095 9399 28101
rect 9858 28092 9864 28104
rect 9916 28092 9922 28144
rect 10229 28135 10287 28141
rect 10229 28101 10241 28135
rect 10275 28132 10287 28135
rect 10502 28132 10508 28144
rect 10275 28104 10508 28132
rect 10275 28101 10287 28104
rect 10229 28095 10287 28101
rect 10502 28092 10508 28104
rect 10560 28092 10566 28144
rect 5776 28036 5821 28064
rect 7668 28036 8248 28064
rect 8481 28067 8539 28073
rect 5776 28024 5782 28036
rect 8481 28033 8493 28067
rect 8527 28033 8539 28067
rect 8481 28027 8539 28033
rect 8665 28067 8723 28073
rect 8665 28033 8677 28067
rect 8711 28064 8723 28067
rect 10045 28067 10103 28073
rect 8711 28036 9444 28064
rect 8711 28033 8723 28036
rect 8665 28027 8723 28033
rect 1578 27956 1584 28008
rect 1636 27996 1642 28008
rect 2130 27996 2136 28008
rect 1636 27968 2136 27996
rect 1636 27956 1642 27968
rect 2130 27956 2136 27968
rect 2188 27956 2194 28008
rect 4798 27996 4804 28008
rect 4759 27968 4804 27996
rect 4798 27956 4804 27968
rect 4856 27956 4862 28008
rect 4893 27999 4951 28005
rect 4893 27965 4905 27999
rect 4939 27965 4951 27999
rect 5166 27996 5172 28008
rect 5127 27968 5172 27996
rect 4893 27959 4951 27965
rect 4065 27931 4123 27937
rect 4065 27897 4077 27931
rect 4111 27928 4123 27931
rect 4706 27928 4712 27940
rect 4111 27900 4712 27928
rect 4111 27897 4123 27900
rect 4065 27891 4123 27897
rect 4706 27888 4712 27900
rect 4764 27888 4770 27940
rect 4908 27928 4936 27959
rect 5166 27956 5172 27968
rect 5224 27956 5230 28008
rect 8202 27956 8208 28008
rect 8260 27996 8266 28008
rect 8496 27996 8524 28027
rect 9416 28008 9444 28036
rect 10045 28033 10057 28067
rect 10091 28064 10103 28067
rect 10410 28064 10416 28076
rect 10091 28036 10416 28064
rect 10091 28033 10103 28036
rect 10045 28027 10103 28033
rect 10410 28024 10416 28036
rect 10468 28064 10474 28076
rect 10962 28064 10968 28076
rect 10468 28036 10968 28064
rect 10468 28024 10474 28036
rect 10962 28024 10968 28036
rect 11020 28024 11026 28076
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 12406 28064 12434 28172
rect 18690 28160 18696 28172
rect 18748 28160 18754 28212
rect 18966 28200 18972 28212
rect 18927 28172 18972 28200
rect 18966 28160 18972 28172
rect 19024 28160 19030 28212
rect 22186 28160 22192 28212
rect 22244 28200 22250 28212
rect 22373 28203 22431 28209
rect 22373 28200 22385 28203
rect 22244 28172 22385 28200
rect 22244 28160 22250 28172
rect 22373 28169 22385 28172
rect 22419 28169 22431 28203
rect 22373 28163 22431 28169
rect 13532 28135 13590 28141
rect 13532 28101 13544 28135
rect 13578 28132 13590 28135
rect 14734 28132 14740 28144
rect 13578 28104 14740 28132
rect 13578 28101 13590 28104
rect 13532 28095 13590 28101
rect 14734 28092 14740 28104
rect 14792 28092 14798 28144
rect 20990 28132 20996 28144
rect 20456 28104 20996 28132
rect 11931 28036 12434 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 12894 28024 12900 28076
rect 12952 28064 12958 28076
rect 13265 28067 13323 28073
rect 13265 28064 13277 28067
rect 12952 28036 13277 28064
rect 12952 28024 12958 28036
rect 13265 28033 13277 28036
rect 13311 28064 13323 28067
rect 14090 28064 14096 28076
rect 13311 28036 14096 28064
rect 13311 28033 13323 28036
rect 13265 28027 13323 28033
rect 14090 28024 14096 28036
rect 14148 28024 14154 28076
rect 16850 28064 16856 28076
rect 16811 28036 16856 28064
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 17126 28064 17132 28076
rect 17087 28036 17132 28064
rect 17126 28024 17132 28036
rect 17184 28024 17190 28076
rect 17773 28067 17831 28073
rect 17773 28033 17785 28067
rect 17819 28064 17831 28067
rect 18138 28064 18144 28076
rect 17819 28036 18144 28064
rect 17819 28033 17831 28036
rect 17773 28027 17831 28033
rect 18138 28024 18144 28036
rect 18196 28064 18202 28076
rect 18509 28067 18567 28073
rect 18509 28064 18521 28067
rect 18196 28036 18521 28064
rect 18196 28024 18202 28036
rect 18509 28033 18521 28036
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 20456 28073 20484 28104
rect 20990 28092 20996 28104
rect 21048 28092 21054 28144
rect 21269 28135 21327 28141
rect 21269 28132 21281 28135
rect 21100 28104 21281 28132
rect 19521 28067 19579 28073
rect 19521 28064 19533 28067
rect 19392 28036 19533 28064
rect 19392 28024 19398 28036
rect 19521 28033 19533 28036
rect 19567 28033 19579 28067
rect 19521 28027 19579 28033
rect 20441 28067 20499 28073
rect 20441 28033 20453 28067
rect 20487 28033 20499 28067
rect 20441 28027 20499 28033
rect 20530 28024 20536 28076
rect 20588 28064 20594 28076
rect 20625 28067 20683 28073
rect 20625 28064 20637 28067
rect 20588 28036 20637 28064
rect 20588 28024 20594 28036
rect 20625 28033 20637 28036
rect 20671 28033 20683 28067
rect 20625 28027 20683 28033
rect 20717 28067 20775 28073
rect 20717 28033 20729 28067
rect 20763 28064 20775 28067
rect 21100 28064 21128 28104
rect 21269 28101 21281 28104
rect 21315 28132 21327 28135
rect 24029 28135 24087 28141
rect 21315 28104 22140 28132
rect 21315 28101 21327 28104
rect 21269 28095 21327 28101
rect 22112 28076 22140 28104
rect 24029 28101 24041 28135
rect 24075 28132 24087 28135
rect 24857 28135 24915 28141
rect 24857 28132 24869 28135
rect 24075 28104 24869 28132
rect 24075 28101 24087 28104
rect 24029 28095 24087 28101
rect 24857 28101 24869 28104
rect 24903 28101 24915 28135
rect 24857 28095 24915 28101
rect 20763 28036 21128 28064
rect 21177 28067 21235 28073
rect 20763 28033 20775 28036
rect 20717 28027 20775 28033
rect 21177 28033 21189 28067
rect 21223 28064 21235 28067
rect 21450 28064 21456 28076
rect 21223 28036 21456 28064
rect 21223 28033 21235 28036
rect 21177 28027 21235 28033
rect 21450 28024 21456 28036
rect 21508 28024 21514 28076
rect 22094 28064 22100 28076
rect 22055 28036 22100 28064
rect 22094 28024 22100 28036
rect 22152 28024 22158 28076
rect 22189 28067 22247 28073
rect 22189 28033 22201 28067
rect 22235 28064 22247 28067
rect 22738 28064 22744 28076
rect 22235 28036 22744 28064
rect 22235 28033 22247 28036
rect 22189 28027 22247 28033
rect 22738 28024 22744 28036
rect 22796 28024 22802 28076
rect 24210 28064 24216 28076
rect 24171 28036 24216 28064
rect 24210 28024 24216 28036
rect 24268 28024 24274 28076
rect 24302 28024 24308 28076
rect 24360 28064 24366 28076
rect 24765 28067 24823 28073
rect 24360 28036 24453 28064
rect 24360 28024 24366 28036
rect 24765 28033 24777 28067
rect 24811 28033 24823 28067
rect 24765 28027 24823 28033
rect 24949 28067 25007 28073
rect 24949 28033 24961 28067
rect 24995 28033 25007 28067
rect 24949 28027 25007 28033
rect 8260 27968 9352 27996
rect 8260 27956 8266 27968
rect 5258 27928 5264 27940
rect 4908 27900 5264 27928
rect 5258 27888 5264 27900
rect 5316 27888 5322 27940
rect 4617 27863 4675 27869
rect 4617 27829 4629 27863
rect 4663 27860 4675 27863
rect 5442 27860 5448 27872
rect 4663 27832 5448 27860
rect 4663 27829 4675 27832
rect 4617 27823 4675 27829
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 7837 27863 7895 27869
rect 7837 27829 7849 27863
rect 7883 27860 7895 27863
rect 8478 27860 8484 27872
rect 7883 27832 8484 27860
rect 7883 27829 7895 27832
rect 7837 27823 7895 27829
rect 8478 27820 8484 27832
rect 8536 27820 8542 27872
rect 9324 27869 9352 27968
rect 9398 27956 9404 28008
rect 9456 27956 9462 28008
rect 11790 27996 11796 28008
rect 11751 27968 11796 27996
rect 11790 27956 11796 27968
rect 11848 27956 11854 28008
rect 12250 27996 12256 28008
rect 12211 27968 12256 27996
rect 12250 27956 12256 27968
rect 12308 27956 12314 28008
rect 15105 27999 15163 28005
rect 15105 27965 15117 27999
rect 15151 27965 15163 27999
rect 15105 27959 15163 27965
rect 15381 27999 15439 28005
rect 15381 27965 15393 27999
rect 15427 27996 15439 27999
rect 15562 27996 15568 28008
rect 15427 27968 15568 27996
rect 15427 27965 15439 27968
rect 15381 27959 15439 27965
rect 14645 27931 14703 27937
rect 14645 27897 14657 27931
rect 14691 27928 14703 27931
rect 15120 27928 15148 27959
rect 15562 27956 15568 27968
rect 15620 27956 15626 28008
rect 16390 27956 16396 28008
rect 16448 27996 16454 28008
rect 16945 27999 17003 28005
rect 16945 27996 16957 27999
rect 16448 27968 16957 27996
rect 16448 27956 16454 27968
rect 16945 27965 16957 27968
rect 16991 27965 17003 27999
rect 24320 27996 24348 28024
rect 16945 27959 17003 27965
rect 24228 27968 24348 27996
rect 15470 27928 15476 27940
rect 14691 27900 15476 27928
rect 14691 27897 14703 27900
rect 14645 27891 14703 27897
rect 15470 27888 15476 27900
rect 15528 27888 15534 27940
rect 18506 27888 18512 27940
rect 18564 27928 18570 27940
rect 19521 27931 19579 27937
rect 19521 27928 19533 27931
rect 18564 27900 19533 27928
rect 18564 27888 18570 27900
rect 19521 27897 19533 27900
rect 19567 27897 19579 27931
rect 19521 27891 19579 27897
rect 20257 27931 20315 27937
rect 20257 27897 20269 27931
rect 20303 27928 20315 27931
rect 24228 27928 24256 27968
rect 24394 27956 24400 28008
rect 24452 27996 24458 28008
rect 24780 27996 24808 28027
rect 24452 27968 24808 27996
rect 24452 27956 24458 27968
rect 24854 27956 24860 28008
rect 24912 27996 24918 28008
rect 24964 27996 24992 28027
rect 24912 27968 24992 27996
rect 24912 27956 24918 27968
rect 20303 27900 24256 27928
rect 20303 27897 20315 27900
rect 20257 27891 20315 27897
rect 9309 27863 9367 27869
rect 9309 27829 9321 27863
rect 9355 27829 9367 27863
rect 9309 27823 9367 27829
rect 16206 27820 16212 27872
rect 16264 27860 16270 27872
rect 16853 27863 16911 27869
rect 16853 27860 16865 27863
rect 16264 27832 16865 27860
rect 16264 27820 16270 27832
rect 16853 27829 16865 27832
rect 16899 27829 16911 27863
rect 16853 27823 16911 27829
rect 16942 27820 16948 27872
rect 17000 27860 17006 27872
rect 17313 27863 17371 27869
rect 17313 27860 17325 27863
rect 17000 27832 17325 27860
rect 17000 27820 17006 27832
rect 17313 27829 17325 27832
rect 17359 27829 17371 27863
rect 17313 27823 17371 27829
rect 17402 27820 17408 27872
rect 17460 27860 17466 27872
rect 17865 27863 17923 27869
rect 17865 27860 17877 27863
rect 17460 27832 17877 27860
rect 17460 27820 17466 27832
rect 17865 27829 17877 27832
rect 17911 27829 17923 27863
rect 18782 27860 18788 27872
rect 18743 27832 18788 27860
rect 17865 27823 17923 27829
rect 18782 27820 18788 27832
rect 18840 27820 18846 27872
rect 19536 27860 19564 27891
rect 21174 27860 21180 27872
rect 19536 27832 21180 27860
rect 21174 27820 21180 27832
rect 21232 27820 21238 27872
rect 21266 27820 21272 27872
rect 21324 27860 21330 27872
rect 22646 27860 22652 27872
rect 21324 27832 22652 27860
rect 21324 27820 21330 27832
rect 22646 27820 22652 27832
rect 22704 27820 22710 27872
rect 24026 27860 24032 27872
rect 23987 27832 24032 27860
rect 24026 27820 24032 27832
rect 24084 27820 24090 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2406 27616 2412 27668
rect 2464 27656 2470 27668
rect 2501 27659 2559 27665
rect 2501 27656 2513 27659
rect 2464 27628 2513 27656
rect 2464 27616 2470 27628
rect 2501 27625 2513 27628
rect 2547 27625 2559 27659
rect 2501 27619 2559 27625
rect 4157 27659 4215 27665
rect 4157 27625 4169 27659
rect 4203 27656 4215 27659
rect 4798 27656 4804 27668
rect 4203 27628 4804 27656
rect 4203 27625 4215 27628
rect 4157 27619 4215 27625
rect 4798 27616 4804 27628
rect 4856 27616 4862 27668
rect 5353 27659 5411 27665
rect 5353 27625 5365 27659
rect 5399 27625 5411 27659
rect 5353 27619 5411 27625
rect 4614 27548 4620 27600
rect 4672 27588 4678 27600
rect 5368 27588 5396 27619
rect 7834 27616 7840 27668
rect 7892 27656 7898 27668
rect 10502 27656 10508 27668
rect 7892 27628 10508 27656
rect 7892 27616 7898 27628
rect 10502 27616 10508 27628
rect 10560 27616 10566 27668
rect 13541 27659 13599 27665
rect 13541 27625 13553 27659
rect 13587 27656 13599 27659
rect 13630 27656 13636 27668
rect 13587 27628 13636 27656
rect 13587 27625 13599 27628
rect 13541 27619 13599 27625
rect 13630 27616 13636 27628
rect 13688 27616 13694 27668
rect 15933 27659 15991 27665
rect 15933 27625 15945 27659
rect 15979 27656 15991 27659
rect 16574 27656 16580 27668
rect 15979 27628 16580 27656
rect 15979 27625 15991 27628
rect 15933 27619 15991 27625
rect 16574 27616 16580 27628
rect 16632 27616 16638 27668
rect 18233 27659 18291 27665
rect 18233 27625 18245 27659
rect 18279 27656 18291 27659
rect 18506 27656 18512 27668
rect 18279 27628 18512 27656
rect 18279 27625 18291 27628
rect 18233 27619 18291 27625
rect 18506 27616 18512 27628
rect 18564 27616 18570 27668
rect 18690 27616 18696 27668
rect 18748 27656 18754 27668
rect 21266 27656 21272 27668
rect 18748 27628 21272 27656
rect 18748 27616 18754 27628
rect 21266 27616 21272 27628
rect 21324 27616 21330 27668
rect 4672 27560 5396 27588
rect 4672 27548 4678 27560
rect 5626 27548 5632 27600
rect 5684 27588 5690 27600
rect 5721 27591 5779 27597
rect 5721 27588 5733 27591
rect 5684 27560 5733 27588
rect 5684 27548 5690 27560
rect 5721 27557 5733 27560
rect 5767 27557 5779 27591
rect 8294 27588 8300 27600
rect 8255 27560 8300 27588
rect 5721 27551 5779 27557
rect 8294 27548 8300 27560
rect 8352 27548 8358 27600
rect 12253 27591 12311 27597
rect 12253 27557 12265 27591
rect 12299 27588 12311 27591
rect 12342 27588 12348 27600
rect 12299 27560 12348 27588
rect 12299 27557 12311 27560
rect 12253 27551 12311 27557
rect 12342 27548 12348 27560
rect 12400 27548 12406 27600
rect 13725 27591 13783 27597
rect 13725 27557 13737 27591
rect 13771 27588 13783 27591
rect 14550 27588 14556 27600
rect 13771 27560 14556 27588
rect 13771 27557 13783 27560
rect 13725 27551 13783 27557
rect 14550 27548 14556 27560
rect 14608 27548 14614 27600
rect 15010 27588 15016 27600
rect 14752 27560 15016 27588
rect 4890 27520 4896 27532
rect 4356 27492 4896 27520
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27452 1639 27455
rect 1854 27452 1860 27464
rect 1627 27424 1860 27452
rect 1627 27421 1639 27424
rect 1581 27415 1639 27421
rect 1854 27412 1860 27424
rect 1912 27412 1918 27464
rect 2501 27455 2559 27461
rect 2501 27421 2513 27455
rect 2547 27421 2559 27455
rect 2682 27452 2688 27464
rect 2643 27424 2688 27452
rect 2501 27415 2559 27421
rect 2516 27384 2544 27415
rect 2682 27412 2688 27424
rect 2740 27412 2746 27464
rect 4356 27461 4384 27492
rect 4890 27480 4896 27492
rect 4948 27480 4954 27532
rect 7668 27492 8432 27520
rect 4341 27455 4399 27461
rect 4341 27421 4353 27455
rect 4387 27421 4399 27455
rect 4614 27452 4620 27464
rect 4575 27424 4620 27452
rect 4341 27415 4399 27421
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 4801 27455 4859 27461
rect 4801 27421 4813 27455
rect 4847 27452 4859 27455
rect 5074 27452 5080 27464
rect 4847 27424 5080 27452
rect 4847 27421 4859 27424
rect 4801 27415 4859 27421
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 7668 27461 7696 27492
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27421 7711 27455
rect 7834 27452 7840 27464
rect 7795 27424 7840 27452
rect 7653 27415 7711 27421
rect 3970 27384 3976 27396
rect 2516 27356 3976 27384
rect 3970 27344 3976 27356
rect 4028 27344 4034 27396
rect 4982 27344 4988 27396
rect 5040 27384 5046 27396
rect 5276 27384 5304 27415
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 5442 27384 5448 27396
rect 5040 27356 5448 27384
rect 5040 27344 5046 27356
rect 5442 27344 5448 27356
rect 5500 27384 5506 27396
rect 7852 27384 7880 27412
rect 5500 27356 7880 27384
rect 5500 27344 5506 27356
rect 8202 27344 8208 27396
rect 8260 27384 8266 27396
rect 8297 27387 8355 27393
rect 8297 27384 8309 27387
rect 8260 27356 8309 27384
rect 8260 27344 8266 27356
rect 8297 27353 8309 27356
rect 8343 27353 8355 27387
rect 8404 27384 8432 27492
rect 11146 27480 11152 27532
rect 11204 27520 11210 27532
rect 11204 27492 12434 27520
rect 11204 27480 11210 27492
rect 8570 27452 8576 27464
rect 8483 27424 8576 27452
rect 8570 27412 8576 27424
rect 8628 27452 8634 27464
rect 9493 27455 9551 27461
rect 9493 27452 9505 27455
rect 8628 27424 9505 27452
rect 8628 27412 8634 27424
rect 9493 27421 9505 27424
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 11422 27412 11428 27464
rect 11480 27452 11486 27464
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 11480 27424 11529 27452
rect 11480 27412 11486 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 11793 27455 11851 27461
rect 11793 27421 11805 27455
rect 11839 27452 11851 27455
rect 11974 27452 11980 27464
rect 11839 27424 11980 27452
rect 11839 27421 11851 27424
rect 11793 27415 11851 27421
rect 11974 27412 11980 27424
rect 12032 27412 12038 27464
rect 9125 27387 9183 27393
rect 9125 27384 9137 27387
rect 8404 27356 9137 27384
rect 8297 27347 8355 27353
rect 9125 27353 9137 27356
rect 9171 27384 9183 27387
rect 9214 27384 9220 27396
rect 9171 27356 9220 27384
rect 9171 27353 9183 27356
rect 9125 27347 9183 27353
rect 9214 27344 9220 27356
rect 9272 27344 9278 27396
rect 9306 27344 9312 27396
rect 9364 27384 9370 27396
rect 9364 27356 9409 27384
rect 9364 27344 9370 27356
rect 9858 27344 9864 27396
rect 9916 27384 9922 27396
rect 10413 27387 10471 27393
rect 10413 27384 10425 27387
rect 9916 27356 10425 27384
rect 9916 27344 9922 27356
rect 10413 27353 10425 27356
rect 10459 27353 10471 27387
rect 12250 27384 12256 27396
rect 12211 27356 12256 27384
rect 10413 27347 10471 27353
rect 12250 27344 12256 27356
rect 12308 27344 12314 27396
rect 12406 27384 12434 27492
rect 12710 27480 12716 27532
rect 12768 27520 12774 27532
rect 12768 27492 13584 27520
rect 12768 27480 12774 27492
rect 12529 27455 12587 27461
rect 12529 27421 12541 27455
rect 12575 27452 12587 27455
rect 13078 27452 13084 27464
rect 12575 27424 13084 27452
rect 12575 27421 12587 27424
rect 12529 27415 12587 27421
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 13556 27452 13584 27492
rect 13630 27480 13636 27532
rect 13688 27520 13694 27532
rect 14752 27529 14780 27560
rect 15010 27548 15016 27560
rect 15068 27548 15074 27600
rect 15194 27548 15200 27600
rect 15252 27588 15258 27600
rect 16117 27591 16175 27597
rect 16117 27588 16129 27591
rect 15252 27560 16129 27588
rect 15252 27548 15258 27560
rect 16117 27557 16129 27560
rect 16163 27557 16175 27591
rect 16117 27551 16175 27557
rect 16206 27548 16212 27600
rect 16264 27588 16270 27600
rect 16761 27591 16819 27597
rect 16761 27588 16773 27591
rect 16264 27560 16773 27588
rect 16264 27548 16270 27560
rect 16761 27557 16773 27560
rect 16807 27588 16819 27591
rect 18598 27588 18604 27600
rect 16807 27560 18604 27588
rect 16807 27557 16819 27560
rect 16761 27551 16819 27557
rect 18598 27548 18604 27560
rect 18656 27548 18662 27600
rect 19426 27588 19432 27600
rect 19306 27560 19432 27588
rect 14461 27523 14519 27529
rect 14461 27520 14473 27523
rect 13688 27492 14473 27520
rect 13688 27480 13694 27492
rect 14461 27489 14473 27492
rect 14507 27489 14519 27523
rect 14461 27483 14519 27489
rect 14737 27523 14795 27529
rect 14737 27489 14749 27523
rect 14783 27489 14795 27523
rect 15562 27520 15568 27532
rect 14737 27483 14795 27489
rect 15120 27492 15568 27520
rect 13722 27452 13728 27464
rect 13556 27424 13728 27452
rect 13722 27412 13728 27424
rect 13780 27412 13786 27464
rect 14274 27412 14280 27464
rect 14332 27452 14338 27464
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 14332 27424 14657 27452
rect 14332 27412 14338 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 14826 27452 14832 27464
rect 14787 27424 14832 27452
rect 14645 27415 14703 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27452 14979 27455
rect 15010 27452 15016 27464
rect 14967 27424 15016 27452
rect 14967 27421 14979 27424
rect 14921 27415 14979 27421
rect 13357 27387 13415 27393
rect 13357 27384 13369 27387
rect 12406 27356 13369 27384
rect 13357 27353 13369 27356
rect 13403 27384 13415 27387
rect 13906 27384 13912 27396
rect 13403 27356 13912 27384
rect 13403 27353 13415 27356
rect 13357 27347 13415 27353
rect 13906 27344 13912 27356
rect 13964 27384 13970 27396
rect 14936 27384 14964 27415
rect 15010 27412 15016 27424
rect 15068 27452 15074 27464
rect 15120 27452 15148 27492
rect 15562 27480 15568 27492
rect 15620 27480 15626 27532
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27520 15899 27523
rect 17034 27520 17040 27532
rect 15887 27492 17040 27520
rect 15887 27489 15899 27492
rect 15841 27483 15899 27489
rect 17034 27480 17040 27492
rect 17092 27480 17098 27532
rect 17218 27520 17224 27532
rect 17179 27492 17224 27520
rect 17218 27480 17224 27492
rect 17276 27480 17282 27532
rect 19306 27520 19334 27560
rect 19426 27548 19432 27560
rect 19484 27588 19490 27600
rect 19705 27591 19763 27597
rect 19705 27588 19717 27591
rect 19484 27560 19717 27588
rect 19484 27548 19490 27560
rect 19705 27557 19717 27560
rect 19751 27588 19763 27591
rect 20530 27588 20536 27600
rect 19751 27560 20536 27588
rect 19751 27557 19763 27560
rect 19705 27551 19763 27557
rect 20530 27548 20536 27560
rect 20588 27548 20594 27600
rect 20714 27588 20720 27600
rect 20675 27560 20720 27588
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 25130 27588 25136 27600
rect 25091 27560 25136 27588
rect 25130 27548 25136 27560
rect 25188 27548 25194 27600
rect 37826 27588 37832 27600
rect 37787 27560 37832 27588
rect 37826 27548 37832 27560
rect 37884 27548 37890 27600
rect 20438 27520 20444 27532
rect 17328 27492 19334 27520
rect 20399 27492 20444 27520
rect 15470 27452 15476 27464
rect 15068 27424 15148 27452
rect 15431 27424 15476 27452
rect 15068 27412 15074 27424
rect 15470 27412 15476 27424
rect 15528 27412 15534 27464
rect 15933 27455 15991 27461
rect 15933 27421 15945 27455
rect 15979 27452 15991 27455
rect 16114 27452 16120 27464
rect 15979 27424 16120 27452
rect 15979 27421 15991 27424
rect 15933 27415 15991 27421
rect 16114 27412 16120 27424
rect 16172 27412 16178 27464
rect 17328 27461 17356 27492
rect 20438 27480 20444 27492
rect 20496 27480 20502 27532
rect 21542 27520 21548 27532
rect 21503 27492 21548 27520
rect 21542 27480 21548 27492
rect 21600 27480 21606 27532
rect 23474 27520 23480 27532
rect 22066 27492 23480 27520
rect 17313 27455 17371 27461
rect 17313 27452 17325 27455
rect 16684 27424 17325 27452
rect 16684 27384 16712 27424
rect 17313 27421 17325 27424
rect 17359 27421 17371 27455
rect 17954 27452 17960 27464
rect 17915 27424 17960 27452
rect 17313 27415 17371 27421
rect 17954 27412 17960 27424
rect 18012 27412 18018 27464
rect 18138 27452 18144 27464
rect 18099 27424 18144 27452
rect 18138 27412 18144 27424
rect 18196 27412 18202 27464
rect 18230 27412 18236 27464
rect 18288 27452 18294 27464
rect 20349 27455 20407 27461
rect 20349 27452 20361 27455
rect 18288 27424 18333 27452
rect 19536 27424 20361 27452
rect 18288 27412 18294 27424
rect 13964 27356 14964 27384
rect 15304 27356 16712 27384
rect 16761 27387 16819 27393
rect 13964 27344 13970 27356
rect 1762 27316 1768 27328
rect 1723 27288 1768 27316
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 7837 27319 7895 27325
rect 7837 27285 7849 27319
rect 7883 27316 7895 27319
rect 8386 27316 8392 27328
rect 7883 27288 8392 27316
rect 7883 27285 7895 27288
rect 7837 27279 7895 27285
rect 8386 27276 8392 27288
rect 8444 27316 8450 27328
rect 8481 27319 8539 27325
rect 8481 27316 8493 27319
rect 8444 27288 8493 27316
rect 8444 27276 8450 27288
rect 8481 27285 8493 27288
rect 8527 27285 8539 27319
rect 10502 27316 10508 27328
rect 10463 27288 10508 27316
rect 8481 27279 8539 27285
rect 10502 27276 10508 27288
rect 10560 27276 10566 27328
rect 11330 27316 11336 27328
rect 11291 27288 11336 27316
rect 11330 27276 11336 27288
rect 11388 27276 11394 27328
rect 11701 27319 11759 27325
rect 11701 27285 11713 27319
rect 11747 27316 11759 27319
rect 12066 27316 12072 27328
rect 11747 27288 12072 27316
rect 11747 27285 11759 27288
rect 11701 27279 11759 27285
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 12434 27276 12440 27328
rect 12492 27316 12498 27328
rect 13567 27319 13625 27325
rect 12492 27288 12537 27316
rect 12492 27276 12498 27288
rect 13567 27285 13579 27319
rect 13613 27316 13625 27319
rect 14274 27316 14280 27328
rect 13613 27288 14280 27316
rect 13613 27285 13625 27288
rect 13567 27279 13625 27285
rect 14274 27276 14280 27288
rect 14332 27276 14338 27328
rect 14550 27276 14556 27328
rect 14608 27316 14614 27328
rect 15304 27316 15332 27356
rect 16761 27353 16773 27387
rect 16807 27384 16819 27387
rect 16942 27384 16948 27396
rect 16807 27356 16948 27384
rect 16807 27353 16819 27356
rect 16761 27347 16819 27353
rect 16942 27344 16948 27356
rect 17000 27344 17006 27396
rect 17497 27387 17555 27393
rect 17497 27384 17509 27387
rect 17052 27356 17509 27384
rect 14608 27288 15332 27316
rect 14608 27276 14614 27288
rect 15378 27276 15384 27328
rect 15436 27316 15442 27328
rect 17052 27316 17080 27356
rect 17497 27353 17509 27356
rect 17543 27353 17555 27387
rect 17497 27347 17555 27353
rect 17586 27344 17592 27396
rect 17644 27384 17650 27396
rect 17644 27356 18552 27384
rect 17644 27344 17650 27356
rect 15436 27288 17080 27316
rect 15436 27276 15442 27288
rect 17126 27276 17132 27328
rect 17184 27316 17190 27328
rect 18230 27316 18236 27328
rect 17184 27288 18236 27316
rect 17184 27276 17190 27288
rect 18230 27276 18236 27288
rect 18288 27276 18294 27328
rect 18414 27316 18420 27328
rect 18375 27288 18420 27316
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 18524 27316 18552 27356
rect 19334 27344 19340 27396
rect 19392 27384 19398 27396
rect 19536 27393 19564 27424
rect 20349 27421 20361 27424
rect 20395 27421 20407 27455
rect 20349 27415 20407 27421
rect 21637 27455 21695 27461
rect 21637 27421 21649 27455
rect 21683 27452 21695 27455
rect 22066 27452 22094 27492
rect 23474 27480 23480 27492
rect 23532 27480 23538 27532
rect 24857 27523 24915 27529
rect 24857 27489 24869 27523
rect 24903 27520 24915 27523
rect 25038 27520 25044 27532
rect 24903 27492 25044 27520
rect 24903 27489 24915 27492
rect 24857 27483 24915 27489
rect 25038 27480 25044 27492
rect 25096 27480 25102 27532
rect 21683 27424 22094 27452
rect 21683 27421 21695 27424
rect 21637 27415 21695 27421
rect 22646 27412 22652 27464
rect 22704 27452 22710 27464
rect 23385 27455 23443 27461
rect 23385 27452 23397 27455
rect 22704 27424 23397 27452
rect 22704 27412 22710 27424
rect 23385 27421 23397 27424
rect 23431 27421 23443 27455
rect 23385 27415 23443 27421
rect 24026 27412 24032 27464
rect 24084 27452 24090 27464
rect 24765 27455 24823 27461
rect 24765 27452 24777 27455
rect 24084 27424 24777 27452
rect 24084 27412 24090 27424
rect 24765 27421 24777 27424
rect 24811 27421 24823 27455
rect 38010 27452 38016 27464
rect 37971 27424 38016 27452
rect 24765 27415 24823 27421
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 19521 27387 19579 27393
rect 19521 27384 19533 27387
rect 19392 27356 19533 27384
rect 19392 27344 19398 27356
rect 19521 27353 19533 27356
rect 19567 27353 19579 27387
rect 19521 27347 19579 27353
rect 23477 27387 23535 27393
rect 23477 27353 23489 27387
rect 23523 27384 23535 27387
rect 24854 27384 24860 27396
rect 23523 27356 24860 27384
rect 23523 27353 23535 27356
rect 23477 27347 23535 27353
rect 24854 27344 24860 27356
rect 24912 27344 24918 27396
rect 20990 27316 20996 27328
rect 18524 27288 20996 27316
rect 20990 27276 20996 27288
rect 21048 27276 21054 27328
rect 22005 27319 22063 27325
rect 22005 27285 22017 27319
rect 22051 27316 22063 27319
rect 22094 27316 22100 27328
rect 22051 27288 22100 27316
rect 22051 27285 22063 27288
rect 22005 27279 22063 27285
rect 22094 27276 22100 27288
rect 22152 27276 22158 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1854 27112 1860 27124
rect 1815 27084 1860 27112
rect 1854 27072 1860 27084
rect 1912 27072 1918 27124
rect 5350 27112 5356 27124
rect 4080 27084 5356 27112
rect 4080 27053 4108 27084
rect 5350 27072 5356 27084
rect 5408 27072 5414 27124
rect 7834 27072 7840 27124
rect 7892 27112 7898 27124
rect 9306 27112 9312 27124
rect 7892 27084 9312 27112
rect 7892 27072 7898 27084
rect 9306 27072 9312 27084
rect 9364 27112 9370 27124
rect 11149 27115 11207 27121
rect 11149 27112 11161 27115
rect 9364 27084 11161 27112
rect 9364 27072 9370 27084
rect 11149 27081 11161 27084
rect 11195 27081 11207 27115
rect 11974 27112 11980 27124
rect 11935 27084 11980 27112
rect 11149 27075 11207 27081
rect 11974 27072 11980 27084
rect 12032 27072 12038 27124
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 13725 27115 13783 27121
rect 13725 27112 13737 27115
rect 12124 27084 13737 27112
rect 12124 27072 12130 27084
rect 13725 27081 13737 27084
rect 13771 27081 13783 27115
rect 14274 27112 14280 27124
rect 14235 27084 14280 27112
rect 13725 27075 13783 27081
rect 14274 27072 14280 27084
rect 14332 27072 14338 27124
rect 14384 27084 14596 27112
rect 3329 27047 3387 27053
rect 3329 27013 3341 27047
rect 3375 27044 3387 27047
rect 4065 27047 4123 27053
rect 3375 27016 4016 27044
rect 3375 27013 3387 27016
rect 3329 27007 3387 27013
rect 2038 26976 2044 26988
rect 1999 26948 2044 26976
rect 2038 26936 2044 26948
rect 2096 26936 2102 26988
rect 3510 26976 3516 26988
rect 3471 26948 3516 26976
rect 3510 26936 3516 26948
rect 3568 26936 3574 26988
rect 3602 26936 3608 26988
rect 3660 26976 3666 26988
rect 3988 26976 4016 27016
rect 4065 27013 4077 27047
rect 4111 27013 4123 27047
rect 4065 27007 4123 27013
rect 4281 27047 4339 27053
rect 4281 27013 4293 27047
rect 4327 27044 4339 27047
rect 4706 27044 4712 27056
rect 4327 27016 4712 27044
rect 4327 27013 4339 27016
rect 4281 27007 4339 27013
rect 4706 27004 4712 27016
rect 4764 27004 4770 27056
rect 5166 27044 5172 27056
rect 5079 27016 5172 27044
rect 4982 26976 4988 26988
rect 3660 26948 3705 26976
rect 3988 26948 4988 26976
rect 3660 26936 3666 26948
rect 4982 26936 4988 26948
rect 5040 26936 5046 26988
rect 5092 26985 5120 27016
rect 5166 27004 5172 27016
rect 5224 27044 5230 27056
rect 5534 27044 5540 27056
rect 5224 27016 5540 27044
rect 5224 27004 5230 27016
rect 5534 27004 5540 27016
rect 5592 27004 5598 27056
rect 6454 27044 6460 27056
rect 6012 27016 6460 27044
rect 5077 26979 5135 26985
rect 5077 26945 5089 26979
rect 5123 26945 5135 26979
rect 5258 26976 5264 26988
rect 5219 26948 5264 26976
rect 5077 26939 5135 26945
rect 5258 26936 5264 26948
rect 5316 26936 5322 26988
rect 5350 26936 5356 26988
rect 5408 26976 5414 26988
rect 5810 26976 5816 26988
rect 5408 26948 5453 26976
rect 5771 26948 5816 26976
rect 5408 26936 5414 26948
rect 5810 26936 5816 26948
rect 5868 26936 5874 26988
rect 6012 26985 6040 27016
rect 6454 27004 6460 27016
rect 6512 27044 6518 27056
rect 10036 27047 10094 27053
rect 6512 27016 8248 27044
rect 6512 27004 6518 27016
rect 8220 26988 8248 27016
rect 10036 27013 10048 27047
rect 10082 27044 10094 27047
rect 11330 27044 11336 27056
rect 10082 27016 11336 27044
rect 10082 27013 10094 27016
rect 10036 27007 10094 27013
rect 11330 27004 11336 27016
rect 11388 27004 11394 27056
rect 12345 27047 12403 27053
rect 12345 27013 12357 27047
rect 12391 27044 12403 27047
rect 12710 27044 12716 27056
rect 12391 27016 12716 27044
rect 12391 27013 12403 27016
rect 12345 27007 12403 27013
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 13173 27047 13231 27053
rect 13173 27013 13185 27047
rect 13219 27044 13231 27047
rect 13906 27044 13912 27056
rect 13219 27016 13912 27044
rect 13219 27013 13231 27016
rect 13173 27007 13231 27013
rect 13906 27004 13912 27016
rect 13964 27004 13970 27056
rect 5997 26979 6055 26985
rect 5997 26945 6009 26979
rect 6043 26945 6055 26979
rect 5997 26939 6055 26945
rect 6178 26936 6184 26988
rect 6236 26976 6242 26988
rect 6805 26979 6863 26985
rect 6805 26976 6817 26979
rect 6236 26948 6817 26976
rect 6236 26936 6242 26948
rect 6805 26945 6817 26948
rect 6851 26945 6863 26979
rect 6805 26939 6863 26945
rect 8202 26936 8208 26988
rect 8260 26976 8266 26988
rect 8260 26948 8708 26976
rect 8260 26936 8266 26948
rect 8680 26920 8708 26948
rect 9398 26936 9404 26988
rect 9456 26976 9462 26988
rect 12161 26979 12219 26985
rect 12161 26976 12173 26979
rect 9456 26948 12173 26976
rect 9456 26936 9462 26948
rect 12161 26945 12173 26948
rect 12207 26945 12219 26979
rect 12161 26939 12219 26945
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26945 12495 26979
rect 12437 26939 12495 26945
rect 12897 26979 12955 26985
rect 12897 26945 12909 26979
rect 12943 26976 12955 26979
rect 13630 26976 13636 26988
rect 12943 26948 13492 26976
rect 13591 26948 13636 26976
rect 12943 26945 12955 26948
rect 12897 26939 12955 26945
rect 3878 26868 3884 26920
rect 3936 26908 3942 26920
rect 6549 26911 6607 26917
rect 6549 26908 6561 26911
rect 3936 26880 6561 26908
rect 3936 26868 3942 26880
rect 6549 26877 6561 26880
rect 6595 26877 6607 26911
rect 8389 26911 8447 26917
rect 8389 26908 8401 26911
rect 6549 26871 6607 26877
rect 7944 26880 8401 26908
rect 4798 26840 4804 26852
rect 4264 26812 4804 26840
rect 3326 26772 3332 26784
rect 3287 26744 3332 26772
rect 3326 26732 3332 26744
rect 3384 26732 3390 26784
rect 4264 26781 4292 26812
rect 4798 26800 4804 26812
rect 4856 26800 4862 26852
rect 7742 26800 7748 26852
rect 7800 26840 7806 26852
rect 7944 26849 7972 26880
rect 8389 26877 8401 26880
rect 8435 26877 8447 26911
rect 8662 26908 8668 26920
rect 8575 26880 8668 26908
rect 8389 26871 8447 26877
rect 8662 26868 8668 26880
rect 8720 26908 8726 26920
rect 9582 26908 9588 26920
rect 8720 26880 9588 26908
rect 8720 26868 8726 26880
rect 9582 26868 9588 26880
rect 9640 26868 9646 26920
rect 9674 26868 9680 26920
rect 9732 26908 9738 26920
rect 9769 26911 9827 26917
rect 9769 26908 9781 26911
rect 9732 26880 9781 26908
rect 9732 26868 9738 26880
rect 9769 26877 9781 26880
rect 9815 26877 9827 26911
rect 9769 26871 9827 26877
rect 7929 26843 7987 26849
rect 7929 26840 7941 26843
rect 7800 26812 7941 26840
rect 7800 26800 7806 26812
rect 7929 26809 7941 26812
rect 7975 26809 7987 26843
rect 7929 26803 7987 26809
rect 4249 26775 4307 26781
rect 4249 26741 4261 26775
rect 4295 26741 4307 26775
rect 4249 26735 4307 26741
rect 4433 26775 4491 26781
rect 4433 26741 4445 26775
rect 4479 26772 4491 26775
rect 4614 26772 4620 26784
rect 4479 26744 4620 26772
rect 4479 26741 4491 26744
rect 4433 26735 4491 26741
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 4890 26772 4896 26784
rect 4851 26744 4896 26772
rect 4890 26732 4896 26744
rect 4948 26732 4954 26784
rect 5902 26772 5908 26784
rect 5863 26744 5908 26772
rect 5902 26732 5908 26744
rect 5960 26732 5966 26784
rect 12452 26772 12480 26939
rect 12989 26843 13047 26849
rect 12989 26809 13001 26843
rect 13035 26840 13047 26843
rect 13464 26840 13492 26948
rect 13630 26936 13636 26948
rect 13688 26936 13694 26988
rect 13722 26936 13728 26988
rect 13780 26976 13786 26988
rect 13817 26979 13875 26985
rect 13817 26976 13829 26979
rect 13780 26948 13829 26976
rect 13780 26936 13786 26948
rect 13817 26945 13829 26948
rect 13863 26945 13875 26979
rect 13817 26939 13875 26945
rect 14384 26908 14412 27084
rect 14458 27004 14464 27056
rect 14516 27004 14522 27056
rect 14568 27044 14596 27084
rect 15562 27072 15568 27124
rect 15620 27112 15626 27124
rect 17402 27112 17408 27124
rect 15620 27084 17408 27112
rect 15620 27072 15626 27084
rect 17402 27072 17408 27084
rect 17460 27072 17466 27124
rect 17954 27072 17960 27124
rect 18012 27112 18018 27124
rect 18012 27084 18644 27112
rect 18012 27072 18018 27084
rect 15933 27047 15991 27053
rect 14568 27016 15608 27044
rect 14476 26976 14504 27004
rect 14553 26979 14611 26985
rect 14553 26976 14565 26979
rect 14476 26948 14565 26976
rect 14553 26945 14565 26948
rect 14599 26945 14611 26979
rect 14553 26939 14611 26945
rect 14737 26979 14795 26985
rect 14737 26945 14749 26979
rect 14783 26976 14795 26979
rect 15194 26976 15200 26988
rect 14783 26948 15200 26976
rect 14783 26945 14795 26948
rect 14737 26939 14795 26945
rect 15194 26936 15200 26948
rect 15252 26936 15258 26988
rect 15289 26979 15347 26985
rect 15289 26945 15301 26979
rect 15335 26976 15347 26979
rect 15470 26976 15476 26988
rect 15335 26948 15476 26976
rect 15335 26945 15347 26948
rect 15289 26939 15347 26945
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 15580 26976 15608 27016
rect 15933 27013 15945 27047
rect 15979 27044 15991 27047
rect 18414 27044 18420 27056
rect 15979 27016 18420 27044
rect 15979 27013 15991 27016
rect 15933 27007 15991 27013
rect 18414 27004 18420 27016
rect 18472 27004 18478 27056
rect 18616 27044 18644 27084
rect 19334 27072 19340 27124
rect 19392 27112 19398 27124
rect 20257 27115 20315 27121
rect 20257 27112 20269 27115
rect 19392 27084 20269 27112
rect 19392 27072 19398 27084
rect 20257 27081 20269 27084
rect 20303 27081 20315 27115
rect 20257 27075 20315 27081
rect 20272 27044 20300 27075
rect 24210 27072 24216 27124
rect 24268 27112 24274 27124
rect 24489 27115 24547 27121
rect 24489 27112 24501 27115
rect 24268 27084 24501 27112
rect 24268 27072 24274 27084
rect 24489 27081 24501 27084
rect 24535 27081 24547 27115
rect 24489 27075 24547 27081
rect 20717 27047 20775 27053
rect 20717 27044 20729 27047
rect 18616 27016 20208 27044
rect 20272 27016 20729 27044
rect 16482 26976 16488 26988
rect 15580 26948 16488 26976
rect 16482 26936 16488 26948
rect 16540 26976 16546 26988
rect 16942 26976 16948 26988
rect 16540 26948 16804 26976
rect 16903 26948 16948 26976
rect 16540 26936 16546 26948
rect 14461 26911 14519 26917
rect 14461 26908 14473 26911
rect 14384 26880 14473 26908
rect 14461 26877 14473 26880
rect 14507 26877 14519 26911
rect 14461 26871 14519 26877
rect 14645 26911 14703 26917
rect 14645 26877 14657 26911
rect 14691 26908 14703 26911
rect 15654 26908 15660 26920
rect 14691 26880 15660 26908
rect 14691 26877 14703 26880
rect 14645 26871 14703 26877
rect 15654 26868 15660 26880
rect 15712 26868 15718 26920
rect 16114 26868 16120 26920
rect 16172 26908 16178 26920
rect 16301 26911 16359 26917
rect 16301 26908 16313 26911
rect 16172 26880 16313 26908
rect 16172 26868 16178 26880
rect 16301 26877 16313 26880
rect 16347 26877 16359 26911
rect 16776 26908 16804 26948
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 17589 26979 17647 26985
rect 17589 26945 17601 26979
rect 17635 26976 17647 26979
rect 18230 26976 18236 26988
rect 17635 26948 18236 26976
rect 17635 26945 17647 26948
rect 17589 26939 17647 26945
rect 18230 26936 18236 26948
rect 18288 26936 18294 26988
rect 18966 26936 18972 26988
rect 19024 26976 19030 26988
rect 19133 26979 19191 26985
rect 19133 26976 19145 26979
rect 19024 26948 19145 26976
rect 19024 26936 19030 26948
rect 19133 26945 19145 26948
rect 19179 26945 19191 26979
rect 20180 26976 20208 27016
rect 20717 27013 20729 27016
rect 20763 27013 20775 27047
rect 20917 27047 20975 27053
rect 20917 27044 20929 27047
rect 20717 27007 20775 27013
rect 20824 27016 20929 27044
rect 20824 26976 20852 27016
rect 20917 27013 20929 27016
rect 20963 27013 20975 27047
rect 20917 27007 20975 27013
rect 23661 27047 23719 27053
rect 23661 27013 23673 27047
rect 23707 27044 23719 27047
rect 24946 27044 24952 27056
rect 23707 27016 24952 27044
rect 23707 27013 23719 27016
rect 23661 27007 23719 27013
rect 24946 27004 24952 27016
rect 25004 27004 25010 27056
rect 20180 26948 20852 26976
rect 19133 26939 19191 26945
rect 22094 26936 22100 26988
rect 22152 26976 22158 26988
rect 22281 26979 22339 26985
rect 22152 26948 22197 26976
rect 22152 26936 22158 26948
rect 22281 26945 22293 26979
rect 22327 26945 22339 26979
rect 23842 26976 23848 26988
rect 23803 26948 23848 26976
rect 22281 26939 22339 26945
rect 17865 26911 17923 26917
rect 16776 26880 17816 26908
rect 16301 26871 16359 26877
rect 16209 26843 16267 26849
rect 16209 26840 16221 26843
rect 13035 26812 13400 26840
rect 13464 26812 16221 26840
rect 13035 26809 13047 26812
rect 12989 26803 13047 26809
rect 13081 26775 13139 26781
rect 13081 26772 13093 26775
rect 12452 26744 13093 26772
rect 13081 26741 13093 26744
rect 13127 26772 13139 26775
rect 13262 26772 13268 26784
rect 13127 26744 13268 26772
rect 13127 26741 13139 26744
rect 13081 26735 13139 26741
rect 13262 26732 13268 26744
rect 13320 26732 13326 26784
rect 13372 26772 13400 26812
rect 16209 26809 16221 26812
rect 16255 26840 16267 26843
rect 16390 26840 16396 26852
rect 16255 26812 16396 26840
rect 16255 26809 16267 26812
rect 16209 26803 16267 26809
rect 16390 26800 16396 26812
rect 16448 26800 16454 26852
rect 16850 26840 16856 26852
rect 16592 26812 16856 26840
rect 14826 26772 14832 26784
rect 13372 26744 14832 26772
rect 14826 26732 14832 26744
rect 14884 26732 14890 26784
rect 15381 26775 15439 26781
rect 15381 26741 15393 26775
rect 15427 26772 15439 26775
rect 15470 26772 15476 26784
rect 15427 26744 15476 26772
rect 15427 26741 15439 26744
rect 15381 26735 15439 26741
rect 15470 26732 15476 26744
rect 15528 26732 15534 26784
rect 15930 26772 15936 26784
rect 15891 26744 15936 26772
rect 15930 26732 15936 26744
rect 15988 26732 15994 26784
rect 16114 26732 16120 26784
rect 16172 26772 16178 26784
rect 16592 26772 16620 26812
rect 16850 26800 16856 26812
rect 16908 26840 16914 26852
rect 17678 26840 17684 26852
rect 16908 26812 17684 26840
rect 16908 26800 16914 26812
rect 17678 26800 17684 26812
rect 17736 26800 17742 26852
rect 17788 26840 17816 26880
rect 17865 26877 17877 26911
rect 17911 26908 17923 26911
rect 18138 26908 18144 26920
rect 17911 26880 18144 26908
rect 17911 26877 17923 26880
rect 17865 26871 17923 26877
rect 18138 26868 18144 26880
rect 18196 26908 18202 26920
rect 18874 26908 18880 26920
rect 18196 26880 18552 26908
rect 18835 26880 18880 26908
rect 18196 26868 18202 26880
rect 18414 26840 18420 26852
rect 17788 26812 18420 26840
rect 18414 26800 18420 26812
rect 18472 26800 18478 26852
rect 16172 26744 16620 26772
rect 17037 26775 17095 26781
rect 16172 26732 16178 26744
rect 17037 26741 17049 26775
rect 17083 26772 17095 26775
rect 17494 26772 17500 26784
rect 17083 26744 17500 26772
rect 17083 26741 17095 26744
rect 17037 26735 17095 26741
rect 17494 26732 17500 26744
rect 17552 26732 17558 26784
rect 18524 26772 18552 26880
rect 18874 26868 18880 26880
rect 18932 26868 18938 26920
rect 22296 26852 22324 26939
rect 23842 26936 23848 26948
rect 23900 26936 23906 26988
rect 23937 26979 23995 26985
rect 23937 26945 23949 26979
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 23106 26868 23112 26920
rect 23164 26908 23170 26920
rect 23952 26908 23980 26939
rect 24394 26936 24400 26988
rect 24452 26976 24458 26988
rect 24581 26979 24639 26985
rect 24452 26948 24497 26976
rect 24452 26936 24458 26948
rect 24581 26945 24593 26979
rect 24627 26976 24639 26979
rect 24854 26976 24860 26988
rect 24627 26948 24860 26976
rect 24627 26945 24639 26948
rect 24581 26939 24639 26945
rect 24854 26936 24860 26948
rect 24912 26936 24918 26988
rect 23164 26880 23980 26908
rect 23164 26868 23170 26880
rect 19886 26800 19892 26852
rect 19944 26840 19950 26852
rect 21085 26843 21143 26849
rect 21085 26840 21097 26843
rect 19944 26812 21097 26840
rect 19944 26800 19950 26812
rect 21085 26809 21097 26812
rect 21131 26809 21143 26843
rect 22278 26840 22284 26852
rect 22191 26812 22284 26840
rect 21085 26803 21143 26809
rect 22278 26800 22284 26812
rect 22336 26840 22342 26852
rect 38010 26840 38016 26852
rect 22336 26812 38016 26840
rect 22336 26800 22342 26812
rect 38010 26800 38016 26812
rect 38068 26800 38074 26852
rect 20901 26775 20959 26781
rect 20901 26772 20913 26775
rect 18524 26744 20913 26772
rect 20901 26741 20913 26744
rect 20947 26741 20959 26775
rect 20901 26735 20959 26741
rect 22097 26775 22155 26781
rect 22097 26741 22109 26775
rect 22143 26772 22155 26775
rect 22186 26772 22192 26784
rect 22143 26744 22192 26772
rect 22143 26741 22155 26744
rect 22097 26735 22155 26741
rect 22186 26732 22192 26744
rect 22244 26732 22250 26784
rect 23661 26775 23719 26781
rect 23661 26741 23673 26775
rect 23707 26772 23719 26775
rect 24762 26772 24768 26784
rect 23707 26744 24768 26772
rect 23707 26741 23719 26744
rect 23661 26735 23719 26741
rect 24762 26732 24768 26744
rect 24820 26732 24826 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 3970 26568 3976 26580
rect 3931 26540 3976 26568
rect 3970 26528 3976 26540
rect 4028 26528 4034 26580
rect 5353 26571 5411 26577
rect 5353 26537 5365 26571
rect 5399 26568 5411 26571
rect 5442 26568 5448 26580
rect 5399 26540 5448 26568
rect 5399 26537 5411 26540
rect 5353 26531 5411 26537
rect 5442 26528 5448 26540
rect 5500 26528 5506 26580
rect 6178 26568 6184 26580
rect 6139 26540 6184 26568
rect 6178 26528 6184 26540
rect 6236 26528 6242 26580
rect 9214 26528 9220 26580
rect 9272 26568 9278 26580
rect 10873 26571 10931 26577
rect 10873 26568 10885 26571
rect 9272 26540 10885 26568
rect 9272 26528 9278 26540
rect 10873 26537 10885 26540
rect 10919 26537 10931 26571
rect 12250 26568 12256 26580
rect 12211 26540 12256 26568
rect 10873 26531 10931 26537
rect 3329 26503 3387 26509
rect 3329 26469 3341 26503
rect 3375 26500 3387 26503
rect 3510 26500 3516 26512
rect 3375 26472 3516 26500
rect 3375 26469 3387 26472
rect 3329 26463 3387 26469
rect 3510 26460 3516 26472
rect 3568 26500 3574 26512
rect 5074 26500 5080 26512
rect 3568 26472 5080 26500
rect 3568 26460 3574 26472
rect 5074 26460 5080 26472
rect 5132 26460 5138 26512
rect 5534 26460 5540 26512
rect 5592 26500 5598 26512
rect 8021 26503 8079 26509
rect 8021 26500 8033 26503
rect 5592 26472 8033 26500
rect 5592 26460 5598 26472
rect 8021 26469 8033 26472
rect 8067 26469 8079 26503
rect 8021 26463 8079 26469
rect 4525 26435 4583 26441
rect 4525 26401 4537 26435
rect 4571 26432 4583 26435
rect 5166 26432 5172 26444
rect 4571 26404 5172 26432
rect 4571 26401 4583 26404
rect 4525 26395 4583 26401
rect 5166 26392 5172 26404
rect 5224 26392 5230 26444
rect 5902 26392 5908 26444
rect 5960 26432 5966 26444
rect 7742 26432 7748 26444
rect 5960 26404 6684 26432
rect 7703 26404 7748 26432
rect 5960 26392 5966 26404
rect 1578 26324 1584 26376
rect 1636 26364 1642 26376
rect 1949 26367 2007 26373
rect 1949 26364 1961 26367
rect 1636 26336 1961 26364
rect 1636 26324 1642 26336
rect 1949 26333 1961 26336
rect 1995 26364 2007 26367
rect 3878 26364 3884 26376
rect 1995 26336 3884 26364
rect 1995 26333 2007 26336
rect 1949 26327 2007 26333
rect 3878 26324 3884 26336
rect 3936 26324 3942 26376
rect 4154 26324 4160 26376
rect 4212 26364 4218 26376
rect 4212 26336 4254 26364
rect 4212 26324 4218 26336
rect 4614 26324 4620 26376
rect 4672 26364 4678 26376
rect 5074 26364 5080 26376
rect 4672 26336 4717 26364
rect 5035 26336 5080 26364
rect 4672 26324 4678 26336
rect 5074 26324 5080 26336
rect 5132 26324 5138 26376
rect 6454 26364 6460 26376
rect 6415 26336 6460 26364
rect 6454 26324 6460 26336
rect 6512 26324 6518 26376
rect 6656 26373 6684 26404
rect 7742 26392 7748 26404
rect 7800 26392 7806 26444
rect 7837 26435 7895 26441
rect 7837 26401 7849 26435
rect 7883 26432 7895 26435
rect 8570 26432 8576 26444
rect 7883 26404 8576 26432
rect 7883 26401 7895 26404
rect 7837 26395 7895 26401
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 10888 26432 10916 26531
rect 12250 26528 12256 26540
rect 12308 26528 12314 26580
rect 13078 26568 13084 26580
rect 13039 26540 13084 26568
rect 13078 26528 13084 26540
rect 13136 26528 13142 26580
rect 14550 26528 14556 26580
rect 14608 26528 14614 26580
rect 14737 26571 14795 26577
rect 14737 26537 14749 26571
rect 14783 26537 14795 26571
rect 14918 26568 14924 26580
rect 14879 26540 14924 26568
rect 14737 26531 14795 26537
rect 14568 26500 14596 26528
rect 12406 26472 14596 26500
rect 14752 26500 14780 26531
rect 14918 26528 14924 26540
rect 14976 26528 14982 26580
rect 15562 26568 15568 26580
rect 15028 26540 15568 26568
rect 15028 26500 15056 26540
rect 15562 26528 15568 26540
rect 15620 26528 15626 26580
rect 15838 26528 15844 26580
rect 15896 26568 15902 26580
rect 16209 26571 16267 26577
rect 16209 26568 16221 26571
rect 15896 26540 16221 26568
rect 15896 26528 15902 26540
rect 16209 26537 16221 26540
rect 16255 26537 16267 26571
rect 16209 26531 16267 26537
rect 18046 26528 18052 26580
rect 18104 26568 18110 26580
rect 18322 26568 18328 26580
rect 18104 26540 18149 26568
rect 18283 26540 18328 26568
rect 18104 26528 18110 26540
rect 18322 26528 18328 26540
rect 18380 26528 18386 26580
rect 18874 26528 18880 26580
rect 18932 26568 18938 26580
rect 21269 26571 21327 26577
rect 18932 26540 20576 26568
rect 18932 26528 18938 26540
rect 20548 26512 20576 26540
rect 21269 26537 21281 26571
rect 21315 26568 21327 26571
rect 25038 26568 25044 26580
rect 21315 26540 24716 26568
rect 24999 26540 25044 26568
rect 21315 26537 21327 26540
rect 21269 26531 21327 26537
rect 14752 26472 15056 26500
rect 16393 26503 16451 26509
rect 11793 26435 11851 26441
rect 11793 26432 11805 26435
rect 10888 26404 11805 26432
rect 11793 26401 11805 26404
rect 11839 26401 11851 26435
rect 11793 26395 11851 26401
rect 6549 26367 6607 26373
rect 6549 26333 6561 26367
rect 6595 26333 6607 26367
rect 6549 26327 6607 26333
rect 6641 26367 6699 26373
rect 6641 26333 6653 26367
rect 6687 26333 6699 26367
rect 6822 26364 6828 26376
rect 6783 26336 6828 26364
rect 6641 26327 6699 26333
rect 2216 26299 2274 26305
rect 2216 26265 2228 26299
rect 2262 26296 2274 26299
rect 2590 26296 2596 26308
rect 2262 26268 2596 26296
rect 2262 26265 2274 26268
rect 2216 26259 2274 26265
rect 2590 26256 2596 26268
rect 2648 26256 2654 26308
rect 3602 26256 3608 26308
rect 3660 26296 3666 26308
rect 4430 26296 4436 26308
rect 3660 26268 4436 26296
rect 3660 26256 3666 26268
rect 4172 26237 4200 26268
rect 4430 26256 4436 26268
rect 4488 26256 4494 26308
rect 5718 26256 5724 26308
rect 5776 26296 5782 26308
rect 6564 26296 6592 26327
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 9493 26367 9551 26373
rect 9493 26333 9505 26367
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 7282 26296 7288 26308
rect 5776 26268 7288 26296
rect 5776 26256 5782 26268
rect 7282 26256 7288 26268
rect 7340 26256 7346 26308
rect 7377 26299 7435 26305
rect 7377 26265 7389 26299
rect 7423 26296 7435 26299
rect 8386 26296 8392 26308
rect 7423 26268 8392 26296
rect 7423 26265 7435 26268
rect 7377 26259 7435 26265
rect 8386 26256 8392 26268
rect 8444 26256 8450 26308
rect 9508 26296 9536 26327
rect 9582 26324 9588 26376
rect 9640 26364 9646 26376
rect 11885 26367 11943 26373
rect 9640 26336 9996 26364
rect 9640 26324 9646 26336
rect 9766 26305 9772 26308
rect 8496 26268 9720 26296
rect 4157 26231 4215 26237
rect 4157 26197 4169 26231
rect 4203 26197 4215 26231
rect 4157 26191 4215 26197
rect 5350 26188 5356 26240
rect 5408 26228 5414 26240
rect 5537 26231 5595 26237
rect 5537 26228 5549 26231
rect 5408 26200 5549 26228
rect 5408 26188 5414 26200
rect 5537 26197 5549 26200
rect 5583 26197 5595 26231
rect 5537 26191 5595 26197
rect 8018 26188 8024 26240
rect 8076 26228 8082 26240
rect 8496 26228 8524 26268
rect 9692 26240 9720 26268
rect 9760 26259 9772 26305
rect 9824 26296 9830 26308
rect 9968 26296 9996 26336
rect 11885 26333 11897 26367
rect 11931 26364 11943 26367
rect 12406 26364 12434 26472
rect 14458 26432 14464 26444
rect 13556 26404 14464 26432
rect 13556 26373 13584 26404
rect 14458 26392 14464 26404
rect 14516 26392 14522 26444
rect 11931 26336 12434 26364
rect 13541 26367 13599 26373
rect 11931 26333 11943 26336
rect 11885 26327 11943 26333
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 13722 26364 13728 26376
rect 13683 26336 13728 26364
rect 13541 26327 13599 26333
rect 13722 26324 13728 26336
rect 13780 26324 13786 26376
rect 14568 26364 14596 26472
rect 16393 26469 16405 26503
rect 16439 26469 16451 26503
rect 17034 26500 17040 26512
rect 16995 26472 17040 26500
rect 16393 26463 16451 26469
rect 14645 26435 14703 26441
rect 14645 26401 14657 26435
rect 14691 26432 14703 26435
rect 16114 26432 16120 26444
rect 14691 26404 16120 26432
rect 14691 26401 14703 26404
rect 14645 26395 14703 26401
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 14737 26367 14795 26373
rect 14737 26364 14749 26367
rect 14568 26336 14749 26364
rect 14737 26333 14749 26336
rect 14783 26333 14795 26367
rect 15378 26364 15384 26376
rect 15339 26336 15384 26364
rect 14737 26327 14795 26333
rect 15378 26324 15384 26336
rect 15436 26324 15442 26376
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26333 15623 26367
rect 15565 26327 15623 26333
rect 12066 26296 12072 26308
rect 9824 26268 9860 26296
rect 9968 26268 12072 26296
rect 9766 26256 9772 26259
rect 9824 26256 9830 26268
rect 12066 26256 12072 26268
rect 12124 26296 12130 26308
rect 12713 26299 12771 26305
rect 12713 26296 12725 26299
rect 12124 26268 12725 26296
rect 12124 26256 12130 26268
rect 12713 26265 12725 26268
rect 12759 26265 12771 26299
rect 12894 26296 12900 26308
rect 12855 26268 12900 26296
rect 12713 26259 12771 26265
rect 12894 26256 12900 26268
rect 12952 26296 12958 26308
rect 13446 26296 13452 26308
rect 12952 26268 13452 26296
rect 12952 26256 12958 26268
rect 13446 26256 13452 26268
rect 13504 26256 13510 26308
rect 14461 26299 14519 26305
rect 14461 26265 14473 26299
rect 14507 26265 14519 26299
rect 14461 26259 14519 26265
rect 8076 26200 8524 26228
rect 8076 26188 8082 26200
rect 9674 26188 9680 26240
rect 9732 26188 9738 26240
rect 13725 26231 13783 26237
rect 13725 26197 13737 26231
rect 13771 26228 13783 26231
rect 14476 26228 14504 26259
rect 14550 26256 14556 26308
rect 14608 26296 14614 26308
rect 15580 26296 15608 26327
rect 15930 26324 15936 26376
rect 15988 26364 15994 26376
rect 16408 26364 16436 26463
rect 17034 26460 17040 26472
rect 17092 26460 17098 26512
rect 20530 26460 20536 26512
rect 20588 26500 20594 26512
rect 22094 26500 22100 26512
rect 20588 26472 22100 26500
rect 20588 26460 20594 26472
rect 22094 26460 22100 26472
rect 22152 26460 22158 26512
rect 23474 26500 23480 26512
rect 23435 26472 23480 26500
rect 23474 26460 23480 26472
rect 23532 26460 23538 26512
rect 19334 26432 19340 26444
rect 17788 26404 19340 26432
rect 17788 26373 17816 26404
rect 19334 26392 19340 26404
rect 19392 26392 19398 26444
rect 19797 26435 19855 26441
rect 19797 26432 19809 26435
rect 19444 26404 19809 26432
rect 16853 26367 16911 26373
rect 16853 26364 16865 26367
rect 15988 26336 16160 26364
rect 16408 26336 16865 26364
rect 15988 26324 15994 26336
rect 16022 26296 16028 26308
rect 14608 26268 15608 26296
rect 15983 26268 16028 26296
rect 14608 26256 14614 26268
rect 16022 26256 16028 26268
rect 16080 26256 16086 26308
rect 16132 26296 16160 26336
rect 16853 26333 16865 26336
rect 16899 26333 16911 26367
rect 16853 26327 16911 26333
rect 17681 26367 17739 26373
rect 17681 26333 17693 26367
rect 17727 26333 17739 26367
rect 17681 26327 17739 26333
rect 17773 26367 17831 26373
rect 17773 26333 17785 26367
rect 17819 26333 17831 26367
rect 17773 26327 17831 26333
rect 18141 26367 18199 26373
rect 18141 26333 18153 26367
rect 18187 26364 18199 26367
rect 18230 26364 18236 26376
rect 18187 26336 18236 26364
rect 18187 26333 18199 26336
rect 18141 26327 18199 26333
rect 16225 26299 16283 26305
rect 16225 26296 16237 26299
rect 16132 26268 16237 26296
rect 16225 26265 16237 26268
rect 16271 26265 16283 26299
rect 16225 26259 16283 26265
rect 17310 26256 17316 26308
rect 17368 26296 17374 26308
rect 17696 26296 17724 26327
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 19444 26364 19472 26404
rect 19797 26401 19809 26404
rect 19843 26432 19855 26435
rect 20070 26432 20076 26444
rect 19843 26404 20076 26432
rect 19843 26401 19855 26404
rect 19797 26395 19855 26401
rect 20070 26392 20076 26404
rect 20128 26392 20134 26444
rect 20346 26392 20352 26444
rect 20404 26432 20410 26444
rect 20901 26435 20959 26441
rect 20901 26432 20913 26435
rect 20404 26404 20913 26432
rect 20404 26392 20410 26404
rect 20901 26401 20913 26404
rect 20947 26401 20959 26435
rect 20901 26395 20959 26401
rect 18472 26336 19472 26364
rect 19521 26367 19579 26373
rect 18472 26324 18478 26336
rect 19521 26333 19533 26367
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26364 19671 26367
rect 19886 26364 19892 26376
rect 19659 26336 19892 26364
rect 19659 26333 19671 26336
rect 19613 26327 19671 26333
rect 19536 26296 19564 26327
rect 19886 26324 19892 26336
rect 19944 26324 19950 26376
rect 20990 26364 20996 26376
rect 20951 26336 20996 26364
rect 20990 26324 20996 26336
rect 21048 26324 21054 26376
rect 22112 26373 22140 26460
rect 24688 26441 24716 26540
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 24673 26435 24731 26441
rect 24673 26401 24685 26435
rect 24719 26401 24731 26435
rect 24673 26395 24731 26401
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26333 22155 26367
rect 22353 26367 22411 26373
rect 22353 26364 22365 26367
rect 22097 26327 22155 26333
rect 22296 26336 22365 26364
rect 17368 26268 19932 26296
rect 17368 26256 17374 26268
rect 13771 26200 14504 26228
rect 15473 26231 15531 26237
rect 13771 26197 13783 26200
rect 13725 26191 13783 26197
rect 15473 26197 15485 26231
rect 15519 26228 15531 26231
rect 19242 26228 19248 26240
rect 15519 26200 19248 26228
rect 15519 26197 15531 26200
rect 15473 26191 15531 26197
rect 19242 26188 19248 26200
rect 19300 26188 19306 26240
rect 19904 26228 19932 26268
rect 22186 26256 22192 26308
rect 22244 26296 22250 26308
rect 22296 26296 22324 26336
rect 22353 26333 22365 26336
rect 22399 26333 22411 26367
rect 24762 26364 24768 26376
rect 24723 26336 24768 26364
rect 22353 26327 22411 26333
rect 24762 26324 24768 26336
rect 24820 26324 24826 26376
rect 37182 26324 37188 26376
rect 37240 26364 37246 26376
rect 37461 26367 37519 26373
rect 37461 26364 37473 26367
rect 37240 26336 37473 26364
rect 37240 26324 37246 26336
rect 37461 26333 37473 26336
rect 37507 26333 37519 26367
rect 37734 26364 37740 26376
rect 37695 26336 37740 26364
rect 37461 26327 37519 26333
rect 37734 26324 37740 26336
rect 37792 26324 37798 26376
rect 22244 26268 22324 26296
rect 22244 26256 22250 26268
rect 21726 26228 21732 26240
rect 19904 26200 21732 26228
rect 21726 26188 21732 26200
rect 21784 26188 21790 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 2590 26024 2596 26036
rect 2551 25996 2596 26024
rect 2590 25984 2596 25996
rect 2648 25984 2654 26036
rect 4249 26027 4307 26033
rect 4249 25993 4261 26027
rect 4295 26024 4307 26027
rect 4614 26024 4620 26036
rect 4295 25996 4620 26024
rect 4295 25993 4307 25996
rect 4249 25987 4307 25993
rect 4614 25984 4620 25996
rect 4672 25984 4678 26036
rect 4798 25984 4804 26036
rect 4856 26024 4862 26036
rect 4909 26027 4967 26033
rect 4909 26024 4921 26027
rect 4856 25996 4921 26024
rect 4856 25984 4862 25996
rect 4909 25993 4921 25996
rect 4955 26024 4967 26027
rect 5629 26027 5687 26033
rect 5629 26024 5641 26027
rect 4955 25996 5641 26024
rect 4955 25993 4967 25996
rect 4909 25987 4967 25993
rect 5629 25993 5641 25996
rect 5675 25993 5687 26027
rect 9858 26024 9864 26036
rect 5629 25987 5687 25993
rect 7668 25996 9864 26024
rect 3326 25956 3332 25968
rect 2516 25928 3332 25956
rect 2516 25897 2544 25928
rect 3326 25916 3332 25928
rect 3384 25916 3390 25968
rect 3881 25959 3939 25965
rect 3881 25925 3893 25959
rect 3927 25956 3939 25959
rect 4522 25956 4528 25968
rect 3927 25928 4528 25956
rect 3927 25925 3939 25928
rect 3881 25919 3939 25925
rect 4522 25916 4528 25928
rect 4580 25916 4586 25968
rect 4709 25959 4767 25965
rect 4709 25925 4721 25959
rect 4755 25956 4767 25959
rect 4755 25928 5212 25956
rect 4755 25925 4767 25928
rect 4709 25919 4767 25925
rect 2501 25891 2559 25897
rect 2501 25857 2513 25891
rect 2547 25857 2559 25891
rect 2682 25888 2688 25900
rect 2643 25860 2688 25888
rect 2501 25851 2559 25857
rect 2682 25848 2688 25860
rect 2740 25848 2746 25900
rect 4062 25888 4068 25900
rect 4023 25860 4068 25888
rect 4062 25848 4068 25860
rect 4120 25848 4126 25900
rect 4982 25712 4988 25764
rect 5040 25752 5046 25764
rect 5077 25755 5135 25761
rect 5077 25752 5089 25755
rect 5040 25724 5089 25752
rect 5040 25712 5046 25724
rect 5077 25721 5089 25724
rect 5123 25721 5135 25755
rect 5184 25752 5212 25928
rect 5258 25916 5264 25968
rect 5316 25956 5322 25968
rect 5316 25928 5856 25956
rect 5316 25916 5322 25928
rect 5534 25888 5540 25900
rect 5495 25860 5540 25888
rect 5534 25848 5540 25860
rect 5592 25848 5598 25900
rect 5828 25897 5856 25928
rect 7668 25900 7696 25996
rect 9858 25984 9864 25996
rect 9916 25984 9922 26036
rect 12253 26027 12311 26033
rect 12253 25993 12265 26027
rect 12299 26024 12311 26027
rect 12434 26024 12440 26036
rect 12299 25996 12440 26024
rect 12299 25993 12311 25996
rect 12253 25987 12311 25993
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 15194 26024 15200 26036
rect 14200 25996 15200 26024
rect 10502 25956 10508 25968
rect 8772 25928 10508 25956
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25857 5779 25891
rect 5721 25851 5779 25857
rect 5813 25891 5871 25897
rect 5813 25857 5825 25891
rect 5859 25857 5871 25891
rect 5813 25851 5871 25857
rect 5350 25780 5356 25832
rect 5408 25820 5414 25832
rect 5736 25820 5764 25851
rect 6454 25848 6460 25900
rect 6512 25888 6518 25900
rect 6549 25891 6607 25897
rect 6549 25888 6561 25891
rect 6512 25860 6561 25888
rect 6512 25848 6518 25860
rect 6549 25857 6561 25860
rect 6595 25857 6607 25891
rect 6730 25888 6736 25900
rect 6691 25860 6736 25888
rect 6549 25851 6607 25857
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25857 6883 25891
rect 6825 25851 6883 25857
rect 5408 25792 5764 25820
rect 5408 25780 5414 25792
rect 6638 25780 6644 25832
rect 6696 25820 6702 25832
rect 6840 25820 6868 25851
rect 7098 25848 7104 25900
rect 7156 25888 7162 25900
rect 7466 25888 7472 25900
rect 7156 25860 7472 25888
rect 7156 25848 7162 25860
rect 7466 25848 7472 25860
rect 7524 25848 7530 25900
rect 7650 25888 7656 25900
rect 7611 25860 7656 25888
rect 7650 25848 7656 25860
rect 7708 25848 7714 25900
rect 8570 25848 8576 25900
rect 8628 25888 8634 25900
rect 8665 25891 8723 25897
rect 8665 25888 8677 25891
rect 8628 25860 8677 25888
rect 8628 25848 8634 25860
rect 8665 25857 8677 25860
rect 8711 25857 8723 25891
rect 8665 25851 8723 25857
rect 8772 25832 8800 25928
rect 10502 25916 10508 25928
rect 10560 25956 10566 25968
rect 10689 25959 10747 25965
rect 10689 25956 10701 25959
rect 10560 25928 10701 25956
rect 10560 25916 10566 25928
rect 10689 25925 10701 25928
rect 10735 25925 10747 25959
rect 10689 25919 10747 25925
rect 8846 25848 8852 25900
rect 8904 25888 8910 25900
rect 9493 25891 9551 25897
rect 9493 25888 9505 25891
rect 8904 25860 9505 25888
rect 8904 25848 8910 25860
rect 9493 25857 9505 25860
rect 9539 25857 9551 25891
rect 9674 25888 9680 25900
rect 9635 25860 9680 25888
rect 9493 25851 9551 25857
rect 9674 25848 9680 25860
rect 9732 25848 9738 25900
rect 9769 25891 9827 25897
rect 9769 25857 9781 25891
rect 9815 25857 9827 25891
rect 12066 25888 12072 25900
rect 12027 25860 12072 25888
rect 9769 25851 9827 25857
rect 8754 25820 8760 25832
rect 6696 25792 6868 25820
rect 8715 25792 8760 25820
rect 6696 25780 6702 25792
rect 8754 25780 8760 25792
rect 8812 25780 8818 25832
rect 9784 25820 9812 25851
rect 12066 25848 12072 25860
rect 12124 25848 12130 25900
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25888 12311 25891
rect 12894 25888 12900 25900
rect 12299 25860 12900 25888
rect 12299 25857 12311 25860
rect 12253 25851 12311 25857
rect 12894 25848 12900 25860
rect 12952 25848 12958 25900
rect 13262 25888 13268 25900
rect 13223 25860 13268 25888
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 13449 25891 13507 25897
rect 13449 25857 13461 25891
rect 13495 25888 13507 25891
rect 13630 25888 13636 25900
rect 13495 25860 13636 25888
rect 13495 25857 13507 25860
rect 13449 25851 13507 25857
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 14200 25897 14228 25996
rect 15194 25984 15200 25996
rect 15252 25984 15258 26036
rect 18966 26024 18972 26036
rect 18927 25996 18972 26024
rect 18966 25984 18972 25996
rect 19024 25984 19030 26036
rect 20438 25984 20444 26036
rect 20496 26024 20502 26036
rect 21085 26027 21143 26033
rect 21085 26024 21097 26027
rect 20496 25996 21097 26024
rect 20496 25984 20502 25996
rect 21085 25993 21097 25996
rect 21131 25993 21143 26027
rect 21085 25987 21143 25993
rect 23842 25984 23848 26036
rect 23900 26024 23906 26036
rect 24029 26027 24087 26033
rect 24029 26024 24041 26027
rect 23900 25996 24041 26024
rect 23900 25984 23906 25996
rect 24029 25993 24041 25996
rect 24075 25993 24087 26027
rect 24946 26024 24952 26036
rect 24907 25996 24952 26024
rect 24029 25987 24087 25993
rect 24946 25984 24952 25996
rect 25004 25984 25010 26036
rect 16022 25956 16028 25968
rect 14384 25928 16028 25956
rect 14384 25897 14412 25928
rect 16022 25916 16028 25928
rect 16080 25916 16086 25968
rect 18138 25916 18144 25968
rect 18196 25956 18202 25968
rect 18233 25959 18291 25965
rect 18233 25956 18245 25959
rect 18196 25928 18245 25956
rect 18196 25916 18202 25928
rect 18233 25925 18245 25928
rect 18279 25925 18291 25959
rect 18233 25919 18291 25925
rect 18417 25959 18475 25965
rect 18417 25925 18429 25959
rect 18463 25956 18475 25959
rect 18598 25956 18604 25968
rect 18463 25928 18604 25956
rect 18463 25925 18475 25928
rect 18417 25919 18475 25925
rect 18598 25916 18604 25928
rect 18656 25916 18662 25968
rect 19242 25956 19248 25968
rect 19203 25928 19248 25956
rect 19242 25916 19248 25928
rect 19300 25916 19306 25968
rect 19475 25959 19533 25965
rect 19475 25925 19487 25959
rect 19521 25956 19533 25959
rect 20162 25956 20168 25968
rect 19521 25928 20168 25956
rect 19521 25925 19533 25928
rect 19475 25919 19533 25925
rect 20162 25916 20168 25928
rect 20220 25916 20226 25968
rect 14185 25891 14243 25897
rect 14185 25857 14197 25891
rect 14231 25857 14243 25891
rect 14185 25851 14243 25857
rect 14369 25891 14427 25897
rect 14369 25857 14381 25891
rect 14415 25857 14427 25891
rect 14826 25888 14832 25900
rect 14787 25860 14832 25888
rect 14369 25851 14427 25857
rect 14826 25848 14832 25860
rect 14884 25848 14890 25900
rect 15010 25888 15016 25900
rect 14971 25860 15016 25888
rect 15010 25848 15016 25860
rect 15068 25848 15074 25900
rect 15746 25888 15752 25900
rect 15707 25860 15752 25888
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25888 17095 25891
rect 17310 25888 17316 25900
rect 17083 25860 17316 25888
rect 17083 25857 17095 25860
rect 17037 25851 17095 25857
rect 17310 25848 17316 25860
rect 17368 25848 17374 25900
rect 19150 25888 19156 25900
rect 19111 25860 19156 25888
rect 19150 25848 19156 25860
rect 19208 25848 19214 25900
rect 19337 25891 19395 25897
rect 19337 25857 19349 25891
rect 19383 25888 19395 25891
rect 19886 25888 19892 25900
rect 19383 25860 19892 25888
rect 19383 25857 19395 25860
rect 19337 25851 19395 25857
rect 19886 25848 19892 25860
rect 19944 25848 19950 25900
rect 20070 25888 20076 25900
rect 20031 25860 20076 25888
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20254 25888 20260 25900
rect 20215 25860 20260 25888
rect 20254 25848 20260 25860
rect 20312 25848 20318 25900
rect 20990 25888 20996 25900
rect 20951 25860 20996 25888
rect 20990 25848 20996 25860
rect 21048 25888 21054 25900
rect 22462 25888 22468 25900
rect 21048 25860 22094 25888
rect 22423 25860 22468 25888
rect 21048 25848 21054 25860
rect 9048 25792 9812 25820
rect 5718 25752 5724 25764
rect 5184 25724 5724 25752
rect 5077 25715 5135 25721
rect 5718 25712 5724 25724
rect 5776 25712 5782 25764
rect 9048 25761 9076 25792
rect 19518 25780 19524 25832
rect 19576 25820 19582 25832
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 19576 25792 19625 25820
rect 19576 25780 19582 25792
rect 19613 25789 19625 25792
rect 19659 25820 19671 25823
rect 19702 25820 19708 25832
rect 19659 25792 19708 25820
rect 19659 25789 19671 25792
rect 19613 25783 19671 25789
rect 19702 25780 19708 25792
rect 19760 25780 19766 25832
rect 19978 25780 19984 25832
rect 20036 25820 20042 25832
rect 20622 25820 20628 25832
rect 20036 25792 20628 25820
rect 20036 25780 20042 25792
rect 20622 25780 20628 25792
rect 20680 25780 20686 25832
rect 22066 25820 22094 25860
rect 22462 25848 22468 25860
rect 22520 25848 22526 25900
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 23569 25891 23627 25897
rect 23569 25888 23581 25891
rect 23532 25860 23581 25888
rect 23532 25848 23538 25860
rect 23569 25857 23581 25860
rect 23615 25888 23627 25891
rect 24394 25888 24400 25900
rect 23615 25860 24400 25888
rect 23615 25857 23627 25860
rect 23569 25851 23627 25857
rect 24394 25848 24400 25860
rect 24452 25888 24458 25900
rect 24489 25891 24547 25897
rect 24489 25888 24501 25891
rect 24452 25860 24501 25888
rect 24452 25848 24458 25860
rect 24489 25857 24501 25860
rect 24535 25857 24547 25891
rect 24489 25851 24547 25857
rect 22738 25820 22744 25832
rect 22066 25792 22744 25820
rect 22738 25780 22744 25792
rect 22796 25820 22802 25832
rect 23290 25820 23296 25832
rect 22796 25792 23296 25820
rect 22796 25780 22802 25792
rect 23290 25780 23296 25792
rect 23348 25780 23354 25832
rect 24670 25820 24676 25832
rect 23400 25792 24676 25820
rect 9033 25755 9091 25761
rect 9033 25721 9045 25755
rect 9079 25721 9091 25755
rect 9033 25715 9091 25721
rect 9493 25755 9551 25761
rect 9493 25721 9505 25755
rect 9539 25752 9551 25755
rect 9766 25752 9772 25764
rect 9539 25724 9772 25752
rect 9539 25721 9551 25724
rect 9493 25715 9551 25721
rect 9766 25712 9772 25724
rect 9824 25712 9830 25764
rect 9858 25712 9864 25764
rect 9916 25752 9922 25764
rect 15933 25755 15991 25761
rect 15933 25752 15945 25755
rect 9916 25724 15945 25752
rect 9916 25712 9922 25724
rect 15933 25721 15945 25724
rect 15979 25752 15991 25755
rect 23400 25752 23428 25792
rect 24670 25780 24676 25792
rect 24728 25780 24734 25832
rect 24765 25755 24823 25761
rect 24765 25752 24777 25755
rect 15979 25724 23428 25752
rect 23768 25724 24777 25752
rect 15979 25721 15991 25724
rect 15933 25715 15991 25721
rect 23768 25696 23796 25724
rect 24765 25721 24777 25724
rect 24811 25721 24823 25755
rect 24765 25715 24823 25721
rect 4890 25684 4896 25696
rect 4851 25656 4896 25684
rect 4890 25644 4896 25656
rect 4948 25644 4954 25696
rect 6549 25687 6607 25693
rect 6549 25653 6561 25687
rect 6595 25684 6607 25687
rect 7006 25684 7012 25696
rect 6595 25656 7012 25684
rect 6595 25653 6607 25656
rect 6549 25647 6607 25653
rect 7006 25644 7012 25656
rect 7064 25644 7070 25696
rect 7558 25644 7564 25696
rect 7616 25684 7622 25696
rect 7837 25687 7895 25693
rect 7837 25684 7849 25687
rect 7616 25656 7849 25684
rect 7616 25644 7622 25656
rect 7837 25653 7849 25656
rect 7883 25653 7895 25687
rect 7837 25647 7895 25653
rect 8294 25644 8300 25696
rect 8352 25684 8358 25696
rect 8665 25687 8723 25693
rect 8665 25684 8677 25687
rect 8352 25656 8677 25684
rect 8352 25644 8358 25656
rect 8665 25653 8677 25656
rect 8711 25653 8723 25687
rect 8665 25647 8723 25653
rect 10042 25644 10048 25696
rect 10100 25684 10106 25696
rect 10781 25687 10839 25693
rect 10781 25684 10793 25687
rect 10100 25656 10793 25684
rect 10100 25644 10106 25656
rect 10781 25653 10793 25656
rect 10827 25653 10839 25687
rect 10781 25647 10839 25653
rect 13170 25644 13176 25696
rect 13228 25684 13234 25696
rect 13265 25687 13323 25693
rect 13265 25684 13277 25687
rect 13228 25656 13277 25684
rect 13228 25644 13234 25656
rect 13265 25653 13277 25656
rect 13311 25653 13323 25687
rect 13630 25684 13636 25696
rect 13591 25656 13636 25684
rect 13265 25647 13323 25653
rect 13630 25644 13636 25656
rect 13688 25644 13694 25696
rect 14277 25687 14335 25693
rect 14277 25653 14289 25687
rect 14323 25684 14335 25687
rect 14366 25684 14372 25696
rect 14323 25656 14372 25684
rect 14323 25653 14335 25656
rect 14277 25647 14335 25653
rect 14366 25644 14372 25656
rect 14424 25644 14430 25696
rect 14642 25644 14648 25696
rect 14700 25684 14706 25696
rect 14829 25687 14887 25693
rect 14829 25684 14841 25687
rect 14700 25656 14841 25684
rect 14700 25644 14706 25656
rect 14829 25653 14841 25656
rect 14875 25653 14887 25687
rect 14829 25647 14887 25653
rect 15197 25687 15255 25693
rect 15197 25653 15209 25687
rect 15243 25684 15255 25687
rect 15286 25684 15292 25696
rect 15243 25656 15292 25684
rect 15243 25653 15255 25656
rect 15197 25647 15255 25653
rect 15286 25644 15292 25656
rect 15344 25644 15350 25696
rect 16850 25644 16856 25696
rect 16908 25684 16914 25696
rect 17129 25687 17187 25693
rect 17129 25684 17141 25687
rect 16908 25656 17141 25684
rect 16908 25644 16914 25656
rect 17129 25653 17141 25656
rect 17175 25653 17187 25687
rect 17129 25647 17187 25653
rect 17497 25687 17555 25693
rect 17497 25653 17509 25687
rect 17543 25684 17555 25687
rect 17678 25684 17684 25696
rect 17543 25656 17684 25684
rect 17543 25653 17555 25656
rect 17497 25647 17555 25653
rect 17678 25644 17684 25656
rect 17736 25644 17742 25696
rect 20070 25684 20076 25696
rect 20031 25656 20076 25684
rect 20070 25644 20076 25656
rect 20128 25644 20134 25696
rect 22646 25684 22652 25696
rect 22607 25656 22652 25684
rect 22646 25644 22652 25656
rect 22704 25644 22710 25696
rect 23750 25684 23756 25696
rect 23711 25656 23756 25684
rect 23750 25644 23756 25656
rect 23808 25644 23814 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 4525 25483 4583 25489
rect 4525 25480 4537 25483
rect 4120 25452 4537 25480
rect 4120 25440 4126 25452
rect 4525 25449 4537 25452
rect 4571 25449 4583 25483
rect 4525 25443 4583 25449
rect 6641 25483 6699 25489
rect 6641 25449 6653 25483
rect 6687 25480 6699 25483
rect 6730 25480 6736 25492
rect 6687 25452 6736 25480
rect 6687 25449 6699 25452
rect 6641 25443 6699 25449
rect 6730 25440 6736 25452
rect 6788 25440 6794 25492
rect 8386 25480 8392 25492
rect 8347 25452 8392 25480
rect 8386 25440 8392 25452
rect 8444 25440 8450 25492
rect 8570 25480 8576 25492
rect 8531 25452 8576 25480
rect 8570 25440 8576 25452
rect 8628 25440 8634 25492
rect 9217 25483 9275 25489
rect 9217 25449 9229 25483
rect 9263 25480 9275 25483
rect 9674 25480 9680 25492
rect 9263 25452 9680 25480
rect 9263 25449 9275 25452
rect 9217 25443 9275 25449
rect 9674 25440 9680 25452
rect 9732 25440 9738 25492
rect 13265 25483 13323 25489
rect 13265 25449 13277 25483
rect 13311 25480 13323 25483
rect 13354 25480 13360 25492
rect 13311 25452 13360 25480
rect 13311 25449 13323 25452
rect 13265 25443 13323 25449
rect 13354 25440 13360 25452
rect 13412 25440 13418 25492
rect 15838 25440 15844 25492
rect 15896 25480 15902 25492
rect 16025 25483 16083 25489
rect 16025 25480 16037 25483
rect 15896 25452 16037 25480
rect 15896 25440 15902 25452
rect 16025 25449 16037 25452
rect 16071 25449 16083 25483
rect 16025 25443 16083 25449
rect 19150 25440 19156 25492
rect 19208 25480 19214 25492
rect 19429 25483 19487 25489
rect 19429 25480 19441 25483
rect 19208 25452 19441 25480
rect 19208 25440 19214 25452
rect 19429 25449 19441 25452
rect 19475 25449 19487 25483
rect 20530 25480 20536 25492
rect 19429 25443 19487 25449
rect 20364 25452 20536 25480
rect 5626 25372 5632 25424
rect 5684 25372 5690 25424
rect 5902 25412 5908 25424
rect 5828 25384 5908 25412
rect 4525 25279 4583 25285
rect 4525 25245 4537 25279
rect 4571 25276 4583 25279
rect 4706 25276 4712 25288
rect 4571 25248 4712 25276
rect 4571 25245 4583 25248
rect 4525 25239 4583 25245
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 4798 25236 4804 25288
rect 4856 25276 4862 25288
rect 5644 25285 5672 25372
rect 5537 25279 5595 25285
rect 4856 25248 4901 25276
rect 5537 25254 5549 25279
rect 4856 25236 4862 25248
rect 5460 25245 5549 25254
rect 5583 25245 5595 25279
rect 5460 25239 5595 25245
rect 5626 25279 5684 25285
rect 5626 25245 5638 25279
rect 5672 25245 5684 25279
rect 5626 25239 5684 25245
rect 5742 25279 5800 25285
rect 5742 25245 5754 25279
rect 5788 25276 5800 25279
rect 5828 25276 5856 25384
rect 5902 25372 5908 25384
rect 5960 25372 5966 25424
rect 6086 25372 6092 25424
rect 6144 25412 6150 25424
rect 9858 25412 9864 25424
rect 6144 25384 9864 25412
rect 6144 25372 6150 25384
rect 9858 25372 9864 25384
rect 9916 25372 9922 25424
rect 16945 25415 17003 25421
rect 16945 25381 16957 25415
rect 16991 25412 17003 25415
rect 17862 25412 17868 25424
rect 16991 25384 17868 25412
rect 16991 25381 17003 25384
rect 16945 25375 17003 25381
rect 17862 25372 17868 25384
rect 17920 25372 17926 25424
rect 18601 25415 18659 25421
rect 18601 25381 18613 25415
rect 18647 25381 18659 25415
rect 18601 25375 18659 25381
rect 16114 25344 16120 25356
rect 14292 25316 16120 25344
rect 5788 25248 5856 25276
rect 5905 25279 5963 25285
rect 5788 25245 5800 25248
rect 5742 25239 5800 25245
rect 5905 25245 5917 25279
rect 5951 25276 5963 25279
rect 6822 25276 6828 25288
rect 5951 25248 6828 25276
rect 5951 25245 5963 25248
rect 5905 25239 5963 25245
rect 5460 25226 5580 25239
rect 6822 25236 6828 25248
rect 6880 25276 6886 25288
rect 7190 25276 7196 25288
rect 6880 25248 7196 25276
rect 6880 25236 6886 25248
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 7558 25276 7564 25288
rect 7519 25248 7564 25276
rect 7558 25236 7564 25248
rect 7616 25236 7622 25288
rect 8662 25276 8668 25288
rect 8220 25248 8668 25276
rect 5350 25208 5356 25220
rect 4724 25180 5356 25208
rect 4724 25149 4752 25180
rect 5350 25168 5356 25180
rect 5408 25168 5414 25220
rect 4709 25143 4767 25149
rect 4709 25109 4721 25143
rect 4755 25109 4767 25143
rect 5258 25140 5264 25152
rect 5219 25112 5264 25140
rect 4709 25103 4767 25109
rect 5258 25100 5264 25112
rect 5316 25100 5322 25152
rect 5460 25140 5488 25226
rect 6454 25208 6460 25220
rect 5828 25180 6460 25208
rect 5828 25140 5856 25180
rect 6454 25168 6460 25180
rect 6512 25168 6518 25220
rect 8220 25217 8248 25248
rect 8662 25236 8668 25248
rect 8720 25236 8726 25288
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 8478 25217 8484 25220
rect 8205 25211 8263 25217
rect 8205 25177 8217 25211
rect 8251 25177 8263 25211
rect 8205 25171 8263 25177
rect 8421 25211 8484 25217
rect 8421 25177 8433 25211
rect 8467 25177 8484 25211
rect 8421 25171 8484 25177
rect 8478 25168 8484 25171
rect 8536 25168 8542 25220
rect 9140 25208 9168 25239
rect 9214 25236 9220 25288
rect 9272 25276 9278 25288
rect 9309 25279 9367 25285
rect 9309 25276 9321 25279
rect 9272 25248 9321 25276
rect 9272 25236 9278 25248
rect 9309 25245 9321 25248
rect 9355 25245 9367 25279
rect 9950 25276 9956 25288
rect 9911 25248 9956 25276
rect 9309 25239 9367 25245
rect 9950 25236 9956 25248
rect 10008 25236 10014 25288
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25276 10195 25279
rect 10502 25276 10508 25288
rect 10183 25248 10508 25276
rect 10183 25245 10195 25248
rect 10137 25239 10195 25245
rect 10502 25236 10508 25248
rect 10560 25236 10566 25288
rect 8680 25180 9168 25208
rect 10597 25211 10655 25217
rect 5460 25112 5856 25140
rect 6086 25100 6092 25152
rect 6144 25140 6150 25152
rect 6638 25140 6644 25152
rect 6696 25149 6702 25152
rect 6696 25143 6715 25149
rect 6144 25112 6644 25140
rect 6144 25100 6150 25112
rect 6638 25100 6644 25112
rect 6703 25109 6715 25143
rect 6696 25103 6715 25109
rect 6825 25143 6883 25149
rect 6825 25109 6837 25143
rect 6871 25140 6883 25143
rect 7098 25140 7104 25152
rect 6871 25112 7104 25140
rect 6871 25109 6883 25112
rect 6825 25103 6883 25109
rect 6696 25100 6702 25103
rect 7098 25100 7104 25112
rect 7156 25100 7162 25152
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 7653 25143 7711 25149
rect 7653 25140 7665 25143
rect 7340 25112 7665 25140
rect 7340 25100 7346 25112
rect 7653 25109 7665 25112
rect 7699 25140 7711 25143
rect 8680 25140 8708 25180
rect 10597 25177 10609 25211
rect 10643 25208 10655 25211
rect 10686 25208 10692 25220
rect 10643 25180 10692 25208
rect 10643 25177 10655 25180
rect 10597 25171 10655 25177
rect 10686 25168 10692 25180
rect 10744 25168 10750 25220
rect 10781 25211 10839 25217
rect 10781 25177 10793 25211
rect 10827 25208 10839 25211
rect 11882 25208 11888 25220
rect 10827 25180 11888 25208
rect 10827 25177 10839 25180
rect 10781 25171 10839 25177
rect 11882 25168 11888 25180
rect 11940 25168 11946 25220
rect 12710 25168 12716 25220
rect 12768 25208 12774 25220
rect 13081 25211 13139 25217
rect 13081 25208 13093 25211
rect 12768 25180 13093 25208
rect 12768 25168 12774 25180
rect 13081 25177 13093 25180
rect 13127 25177 13139 25211
rect 13081 25171 13139 25177
rect 13297 25211 13355 25217
rect 13297 25177 13309 25211
rect 13343 25208 13355 25211
rect 14292 25208 14320 25316
rect 16114 25304 16120 25316
rect 16172 25304 16178 25356
rect 16482 25304 16488 25356
rect 16540 25344 16546 25356
rect 17402 25344 17408 25356
rect 16540 25316 17408 25344
rect 16540 25304 16546 25316
rect 17402 25304 17408 25316
rect 17460 25304 17466 25356
rect 17497 25347 17555 25353
rect 17497 25313 17509 25347
rect 17543 25344 17555 25347
rect 18506 25344 18512 25356
rect 17543 25316 18512 25344
rect 17543 25313 17555 25316
rect 17497 25307 17555 25313
rect 14550 25236 14556 25288
rect 14608 25276 14614 25288
rect 14829 25279 14887 25285
rect 14829 25276 14841 25279
rect 14608 25248 14841 25276
rect 14608 25236 14614 25248
rect 14829 25245 14841 25248
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 15013 25279 15071 25285
rect 15013 25245 15025 25279
rect 15059 25245 15071 25279
rect 15013 25239 15071 25245
rect 13343 25180 14320 25208
rect 13343 25177 13355 25180
rect 13297 25171 13355 25177
rect 14366 25168 14372 25220
rect 14424 25208 14430 25220
rect 15028 25208 15056 25239
rect 16022 25236 16028 25288
rect 16080 25236 16086 25288
rect 17310 25276 17316 25288
rect 17271 25248 17316 25276
rect 17310 25236 17316 25248
rect 17368 25236 17374 25288
rect 14424 25180 15056 25208
rect 15841 25211 15899 25217
rect 14424 25168 14430 25180
rect 15841 25177 15853 25211
rect 15887 25208 15899 25211
rect 16040 25208 16068 25236
rect 17512 25208 17540 25307
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 18616 25344 18644 25375
rect 18874 25372 18880 25424
rect 18932 25412 18938 25424
rect 19334 25412 19340 25424
rect 18932 25384 19340 25412
rect 18932 25372 18938 25384
rect 19334 25372 19340 25384
rect 19392 25372 19398 25424
rect 20364 25353 20392 25452
rect 20530 25440 20536 25452
rect 20588 25440 20594 25492
rect 23014 25440 23020 25492
rect 23072 25480 23078 25492
rect 23109 25483 23167 25489
rect 23109 25480 23121 25483
rect 23072 25452 23121 25480
rect 23072 25440 23078 25452
rect 23109 25449 23121 25452
rect 23155 25449 23167 25483
rect 23109 25443 23167 25449
rect 21726 25412 21732 25424
rect 21639 25384 21732 25412
rect 21726 25372 21732 25384
rect 21784 25412 21790 25424
rect 22462 25412 22468 25424
rect 21784 25384 22468 25412
rect 21784 25372 21790 25384
rect 22462 25372 22468 25384
rect 22520 25412 22526 25424
rect 22520 25384 22784 25412
rect 22520 25372 22526 25384
rect 20349 25347 20407 25353
rect 18616 25316 19478 25344
rect 18874 25276 18880 25288
rect 18835 25248 18880 25276
rect 18874 25236 18880 25248
rect 18932 25236 18938 25288
rect 19450 25285 19478 25316
rect 20349 25313 20361 25347
rect 20395 25313 20407 25347
rect 20349 25307 20407 25313
rect 19429 25279 19487 25285
rect 18984 25248 19380 25276
rect 15887 25180 16068 25208
rect 17328 25180 17540 25208
rect 18601 25211 18659 25217
rect 15887 25177 15899 25180
rect 15841 25171 15899 25177
rect 17328 25152 17356 25180
rect 18601 25177 18613 25211
rect 18647 25208 18659 25211
rect 18984 25208 19012 25248
rect 19352 25220 19380 25248
rect 19429 25245 19441 25279
rect 19475 25245 19487 25279
rect 19429 25239 19487 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25276 19671 25279
rect 19978 25276 19984 25288
rect 19659 25248 19984 25276
rect 19659 25245 19671 25248
rect 19613 25239 19671 25245
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 22756 25285 22784 25384
rect 22830 25304 22836 25356
rect 22888 25344 22894 25356
rect 22888 25316 22933 25344
rect 22888 25304 22894 25316
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25245 22799 25279
rect 22741 25239 22799 25245
rect 18647 25180 19012 25208
rect 18647 25177 18659 25180
rect 18601 25171 18659 25177
rect 19334 25168 19340 25220
rect 19392 25168 19398 25220
rect 19702 25168 19708 25220
rect 19760 25208 19766 25220
rect 20594 25211 20652 25217
rect 20594 25208 20606 25211
rect 19760 25180 20606 25208
rect 19760 25168 19766 25180
rect 20594 25177 20606 25180
rect 20640 25177 20652 25211
rect 20594 25171 20652 25177
rect 10134 25140 10140 25152
rect 7699 25112 8708 25140
rect 10095 25112 10140 25140
rect 7699 25109 7711 25112
rect 7653 25103 7711 25109
rect 10134 25100 10140 25112
rect 10192 25100 10198 25152
rect 10962 25140 10968 25152
rect 10923 25112 10968 25140
rect 10962 25100 10968 25112
rect 11020 25100 11026 25152
rect 13446 25140 13452 25152
rect 13407 25112 13452 25140
rect 13446 25100 13452 25112
rect 13504 25100 13510 25152
rect 14918 25140 14924 25152
rect 14879 25112 14924 25140
rect 14918 25100 14924 25112
rect 14976 25100 14982 25152
rect 15378 25100 15384 25152
rect 15436 25140 15442 25152
rect 16041 25143 16099 25149
rect 16041 25140 16053 25143
rect 15436 25112 16053 25140
rect 15436 25100 15442 25112
rect 16041 25109 16053 25112
rect 16087 25109 16099 25143
rect 16206 25140 16212 25152
rect 16167 25112 16212 25140
rect 16041 25103 16099 25109
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 17310 25100 17316 25152
rect 17368 25100 17374 25152
rect 17954 25100 17960 25152
rect 18012 25140 18018 25152
rect 18690 25140 18696 25152
rect 18012 25112 18696 25140
rect 18012 25100 18018 25112
rect 18690 25100 18696 25112
rect 18748 25140 18754 25152
rect 18785 25143 18843 25149
rect 18785 25140 18797 25143
rect 18748 25112 18797 25140
rect 18748 25100 18754 25112
rect 18785 25109 18797 25112
rect 18831 25109 18843 25143
rect 18785 25103 18843 25109
rect 18874 25100 18880 25152
rect 18932 25140 18938 25152
rect 20714 25140 20720 25152
rect 18932 25112 20720 25140
rect 18932 25100 18938 25112
rect 20714 25100 20720 25112
rect 20772 25100 20778 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 13725 24939 13783 24945
rect 13725 24905 13737 24939
rect 13771 24936 13783 24939
rect 15197 24939 15255 24945
rect 13771 24908 15148 24936
rect 13771 24905 13783 24908
rect 13725 24899 13783 24905
rect 4884 24871 4942 24877
rect 4884 24837 4896 24871
rect 4930 24868 4942 24871
rect 5258 24868 5264 24880
rect 4930 24840 5264 24868
rect 4930 24837 4942 24840
rect 4884 24831 4942 24837
rect 5258 24828 5264 24840
rect 5316 24828 5322 24880
rect 6840 24840 9674 24868
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24800 2283 24803
rect 2314 24800 2320 24812
rect 2271 24772 2320 24800
rect 2271 24769 2283 24772
rect 2225 24763 2283 24769
rect 2314 24760 2320 24772
rect 2372 24760 2378 24812
rect 2406 24760 2412 24812
rect 2464 24800 2470 24812
rect 2682 24800 2688 24812
rect 2464 24772 2688 24800
rect 2464 24760 2470 24772
rect 2682 24760 2688 24772
rect 2740 24760 2746 24812
rect 3142 24800 3148 24812
rect 3103 24772 3148 24800
rect 3142 24760 3148 24772
rect 3200 24760 3206 24812
rect 6454 24760 6460 24812
rect 6512 24800 6518 24812
rect 6840 24809 6868 24840
rect 6825 24803 6883 24809
rect 6825 24800 6837 24803
rect 6512 24772 6837 24800
rect 6512 24760 6518 24772
rect 6825 24769 6837 24772
rect 6871 24769 6883 24803
rect 6825 24763 6883 24769
rect 7926 24760 7932 24812
rect 7984 24800 7990 24812
rect 8277 24803 8335 24809
rect 8277 24800 8289 24803
rect 7984 24772 8289 24800
rect 7984 24760 7990 24772
rect 8277 24769 8289 24772
rect 8323 24769 8335 24803
rect 9646 24800 9674 24840
rect 10134 24828 10140 24880
rect 10192 24868 10198 24880
rect 10413 24871 10471 24877
rect 10413 24868 10425 24871
rect 10192 24840 10425 24868
rect 10192 24828 10198 24840
rect 10413 24837 10425 24840
rect 10459 24837 10471 24871
rect 10413 24831 10471 24837
rect 10505 24871 10563 24877
rect 10505 24837 10517 24871
rect 10551 24868 10563 24871
rect 10962 24868 10968 24880
rect 10551 24840 10968 24868
rect 10551 24837 10563 24840
rect 10505 24831 10563 24837
rect 10962 24828 10968 24840
rect 11020 24828 11026 24880
rect 14366 24868 14372 24880
rect 14327 24840 14372 24868
rect 14366 24828 14372 24840
rect 14424 24828 14430 24880
rect 15120 24868 15148 24908
rect 15197 24905 15209 24939
rect 15243 24936 15255 24939
rect 15746 24936 15752 24948
rect 15243 24908 15752 24936
rect 15243 24905 15255 24908
rect 15197 24899 15255 24905
rect 15746 24896 15752 24908
rect 15804 24896 15810 24948
rect 18874 24936 18880 24948
rect 16868 24908 18880 24936
rect 16868 24868 16896 24908
rect 18874 24896 18880 24908
rect 18932 24896 18938 24948
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19392 24908 19437 24936
rect 19536 24908 20024 24936
rect 19392 24896 19398 24908
rect 17954 24868 17960 24880
rect 15120 24840 16896 24868
rect 17604 24840 17960 24868
rect 9950 24800 9956 24812
rect 9646 24772 9956 24800
rect 8277 24763 8335 24769
rect 9950 24760 9956 24772
rect 10008 24760 10014 24812
rect 10226 24800 10232 24812
rect 10187 24772 10232 24800
rect 10226 24760 10232 24772
rect 10284 24760 10290 24812
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 1578 24692 1584 24744
rect 1636 24732 1642 24744
rect 4617 24735 4675 24741
rect 4617 24732 4629 24735
rect 1636 24704 4629 24732
rect 1636 24692 1642 24704
rect 4617 24701 4629 24704
rect 4663 24701 4675 24735
rect 6549 24735 6607 24741
rect 6549 24732 6561 24735
rect 4617 24695 4675 24701
rect 6012 24704 6561 24732
rect 6012 24676 6040 24704
rect 6549 24701 6561 24704
rect 6595 24701 6607 24735
rect 8018 24732 8024 24744
rect 7979 24704 8024 24732
rect 6549 24695 6607 24701
rect 8018 24692 8024 24704
rect 8076 24692 8082 24744
rect 10042 24732 10048 24744
rect 9048 24704 10048 24732
rect 5994 24664 6000 24676
rect 5907 24636 6000 24664
rect 5994 24624 6000 24636
rect 6052 24624 6058 24676
rect 2222 24596 2228 24608
rect 2183 24568 2228 24596
rect 2222 24556 2228 24568
rect 2280 24556 2286 24608
rect 3050 24556 3056 24608
rect 3108 24596 3114 24608
rect 3237 24599 3295 24605
rect 3237 24596 3249 24599
rect 3108 24568 3249 24596
rect 3108 24556 3114 24568
rect 3237 24565 3249 24568
rect 3283 24565 3295 24599
rect 3602 24596 3608 24608
rect 3563 24568 3608 24596
rect 3237 24559 3295 24565
rect 3602 24556 3608 24568
rect 3660 24556 3666 24608
rect 4890 24556 4896 24608
rect 4948 24596 4954 24608
rect 5258 24596 5264 24608
rect 4948 24568 5264 24596
rect 4948 24556 4954 24568
rect 5258 24556 5264 24568
rect 5316 24596 5322 24608
rect 9048 24596 9076 24704
rect 10042 24692 10048 24704
rect 10100 24692 10106 24744
rect 10612 24732 10640 24763
rect 10686 24760 10692 24812
rect 10744 24800 10750 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 10744 24772 11713 24800
rect 10744 24760 10750 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11882 24800 11888 24812
rect 11843 24772 11888 24800
rect 11701 24763 11759 24769
rect 11882 24760 11888 24772
rect 11940 24760 11946 24812
rect 12710 24760 12716 24812
rect 12768 24800 12774 24812
rect 13449 24803 13507 24809
rect 13449 24800 13461 24803
rect 12768 24772 13461 24800
rect 12768 24760 12774 24772
rect 13449 24769 13461 24772
rect 13495 24769 13507 24803
rect 14550 24800 14556 24812
rect 14511 24772 14556 24800
rect 13449 24763 13507 24769
rect 14550 24760 14556 24772
rect 14608 24760 14614 24812
rect 14734 24800 14740 24812
rect 14695 24772 14740 24800
rect 14734 24760 14740 24772
rect 14792 24760 14798 24812
rect 15378 24800 15384 24812
rect 15339 24772 15384 24800
rect 15378 24760 15384 24772
rect 15436 24760 15442 24812
rect 15657 24803 15715 24809
rect 15657 24769 15669 24803
rect 15703 24800 15715 24803
rect 15841 24803 15899 24809
rect 15703 24772 15792 24800
rect 15703 24769 15715 24772
rect 15657 24763 15715 24769
rect 11793 24735 11851 24741
rect 11793 24732 11805 24735
rect 10612 24704 11805 24732
rect 11793 24701 11805 24704
rect 11839 24701 11851 24735
rect 13265 24735 13323 24741
rect 13265 24732 13277 24735
rect 11793 24695 11851 24701
rect 12406 24704 13277 24732
rect 9766 24624 9772 24676
rect 9824 24664 9830 24676
rect 10686 24664 10692 24676
rect 9824 24636 10692 24664
rect 9824 24624 9830 24636
rect 10686 24624 10692 24636
rect 10744 24664 10750 24676
rect 12406 24664 12434 24704
rect 13265 24701 13277 24704
rect 13311 24732 13323 24735
rect 13354 24732 13360 24744
rect 13311 24704 13360 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 13630 24692 13636 24744
rect 13688 24732 13694 24744
rect 13817 24735 13875 24741
rect 13817 24732 13829 24735
rect 13688 24704 13829 24732
rect 13688 24692 13694 24704
rect 13817 24701 13829 24704
rect 13863 24732 13875 24735
rect 13863 24704 15424 24732
rect 13863 24701 13875 24704
rect 13817 24695 13875 24701
rect 10744 24636 12434 24664
rect 10744 24624 10750 24636
rect 5316 24568 9076 24596
rect 9401 24599 9459 24605
rect 5316 24556 5322 24568
rect 9401 24565 9413 24599
rect 9447 24596 9459 24599
rect 9674 24596 9680 24608
rect 9447 24568 9680 24596
rect 9447 24565 9459 24568
rect 9401 24559 9459 24565
rect 9674 24556 9680 24568
rect 9732 24596 9738 24608
rect 10594 24596 10600 24608
rect 9732 24568 10600 24596
rect 9732 24556 9738 24568
rect 10594 24556 10600 24568
rect 10652 24556 10658 24608
rect 10781 24599 10839 24605
rect 10781 24565 10793 24599
rect 10827 24596 10839 24599
rect 11790 24596 11796 24608
rect 10827 24568 11796 24596
rect 10827 24565 10839 24568
rect 10781 24559 10839 24565
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 15396 24596 15424 24704
rect 15764 24664 15792 24772
rect 15841 24769 15853 24803
rect 15887 24800 15899 24803
rect 16114 24800 16120 24812
rect 15887 24772 16120 24800
rect 15887 24769 15899 24772
rect 15841 24763 15899 24769
rect 16114 24760 16120 24772
rect 16172 24760 16178 24812
rect 17494 24800 17500 24812
rect 17455 24772 17500 24800
rect 17494 24760 17500 24772
rect 17552 24760 17558 24812
rect 17604 24809 17632 24840
rect 17954 24828 17960 24840
rect 18012 24828 18018 24880
rect 18616 24840 19012 24868
rect 17589 24803 17647 24809
rect 17589 24769 17601 24803
rect 17635 24769 17647 24803
rect 17589 24763 17647 24769
rect 17678 24760 17684 24812
rect 17736 24803 17742 24812
rect 17736 24775 17778 24803
rect 17736 24760 17742 24775
rect 17862 24760 17868 24812
rect 17920 24800 17926 24812
rect 18616 24809 18644 24840
rect 18509 24803 18567 24809
rect 17920 24772 17965 24800
rect 17920 24760 17926 24772
rect 18509 24769 18521 24803
rect 18555 24769 18567 24803
rect 18509 24763 18567 24769
rect 18601 24803 18659 24809
rect 18601 24769 18613 24803
rect 18647 24769 18659 24803
rect 18601 24763 18659 24769
rect 18785 24803 18843 24809
rect 18874 24803 18880 24812
rect 18785 24769 18797 24803
rect 18831 24775 18880 24803
rect 18831 24769 18843 24775
rect 18785 24763 18843 24769
rect 17221 24735 17279 24741
rect 17221 24701 17233 24735
rect 17267 24732 17279 24735
rect 18524 24732 18552 24763
rect 18874 24760 18880 24775
rect 18932 24760 18938 24812
rect 17267 24704 18552 24732
rect 18693 24735 18751 24741
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 18693 24701 18705 24735
rect 18739 24732 18751 24735
rect 18984 24732 19012 24840
rect 19242 24760 19248 24812
rect 19300 24800 19306 24812
rect 19536 24809 19564 24908
rect 19823 24871 19881 24877
rect 19823 24868 19835 24871
rect 19812 24837 19835 24868
rect 19869 24837 19881 24871
rect 19996 24868 20024 24908
rect 20254 24896 20260 24948
rect 20312 24936 20318 24948
rect 20533 24939 20591 24945
rect 20533 24936 20545 24939
rect 20312 24908 20545 24936
rect 20312 24896 20318 24908
rect 20533 24905 20545 24908
rect 20579 24905 20591 24939
rect 20533 24899 20591 24905
rect 20714 24896 20720 24948
rect 20772 24936 20778 24948
rect 20772 24908 22784 24936
rect 20772 24896 20778 24908
rect 20070 24868 20076 24880
rect 19996 24840 20076 24868
rect 19812 24834 19881 24837
rect 19521 24803 19579 24809
rect 19300 24772 19478 24800
rect 19300 24760 19306 24772
rect 19334 24732 19340 24744
rect 18739 24704 18920 24732
rect 18984 24704 19340 24732
rect 18739 24701 18751 24704
rect 18693 24695 18751 24701
rect 18325 24667 18383 24673
rect 18325 24664 18337 24667
rect 15764 24636 18337 24664
rect 18325 24633 18337 24636
rect 18371 24633 18383 24667
rect 18782 24664 18788 24676
rect 18325 24627 18383 24633
rect 18708 24636 18788 24664
rect 18708 24596 18736 24636
rect 18782 24624 18788 24636
rect 18840 24624 18846 24676
rect 18892 24664 18920 24704
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 19450 24732 19478 24772
rect 19521 24769 19533 24803
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 19613 24803 19671 24809
rect 19613 24769 19625 24803
rect 19659 24769 19671 24803
rect 19613 24763 19671 24769
rect 19705 24803 19763 24809
rect 19812 24806 19932 24834
rect 20070 24828 20076 24840
rect 20128 24828 20134 24880
rect 22646 24868 22652 24880
rect 21928 24840 22652 24868
rect 19705 24769 19717 24803
rect 19751 24769 19763 24803
rect 19705 24763 19763 24769
rect 19628 24732 19656 24763
rect 19450 24704 19656 24732
rect 19720 24732 19748 24763
rect 19794 24732 19800 24744
rect 19720 24704 19800 24732
rect 19794 24692 19800 24704
rect 19852 24692 19858 24744
rect 19702 24664 19708 24676
rect 18892 24636 19708 24664
rect 19702 24624 19708 24636
rect 19760 24624 19766 24676
rect 19904 24664 19932 24806
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24800 20499 24803
rect 20530 24800 20536 24812
rect 20487 24772 20536 24800
rect 20487 24769 20499 24772
rect 20441 24763 20499 24769
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 20625 24803 20683 24809
rect 20625 24769 20637 24803
rect 20671 24800 20683 24803
rect 21928 24800 21956 24840
rect 22646 24828 22652 24840
rect 22704 24828 22710 24880
rect 22756 24868 22784 24908
rect 22830 24896 22836 24948
rect 22888 24936 22894 24948
rect 23382 24936 23388 24948
rect 22888 24908 23388 24936
rect 22888 24896 22894 24908
rect 23382 24896 23388 24908
rect 23440 24936 23446 24948
rect 23477 24939 23535 24945
rect 23477 24936 23489 24939
rect 23440 24908 23489 24936
rect 23440 24896 23446 24908
rect 23477 24905 23489 24908
rect 23523 24905 23535 24939
rect 23477 24899 23535 24905
rect 24762 24868 24768 24880
rect 22756 24840 24624 24868
rect 24723 24840 24768 24868
rect 24596 24812 24624 24840
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 20671 24772 21956 24800
rect 20671 24769 20683 24772
rect 20625 24763 20683 24769
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 20640 24732 20668 24763
rect 22048 24760 22054 24812
rect 22106 24809 22112 24812
rect 22106 24803 22155 24809
rect 22106 24769 22109 24803
rect 22143 24769 22155 24803
rect 22353 24803 22411 24809
rect 22353 24800 22365 24803
rect 22106 24763 22155 24769
rect 22204 24772 22365 24800
rect 22106 24760 22112 24763
rect 22204 24732 22232 24772
rect 22353 24769 22365 24772
rect 22399 24769 22411 24803
rect 22353 24763 22411 24769
rect 24397 24803 24455 24809
rect 24397 24769 24409 24803
rect 24443 24769 24455 24803
rect 24578 24800 24584 24812
rect 24539 24772 24584 24800
rect 24397 24763 24455 24769
rect 20027 24704 20668 24732
rect 22112 24704 22232 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 22112 24676 22140 24704
rect 20162 24664 20168 24676
rect 19904 24636 20168 24664
rect 20162 24624 20168 24636
rect 20220 24624 20226 24676
rect 22094 24624 22100 24676
rect 22152 24624 22158 24676
rect 24412 24664 24440 24763
rect 24578 24760 24584 24772
rect 24636 24760 24642 24812
rect 23216 24636 24440 24664
rect 15396 24568 18736 24596
rect 19150 24556 19156 24608
rect 19208 24596 19214 24608
rect 23216 24596 23244 24636
rect 19208 24568 23244 24596
rect 19208 24556 19214 24568
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 2314 24352 2320 24404
rect 2372 24392 2378 24404
rect 3973 24395 4031 24401
rect 3973 24392 3985 24395
rect 2372 24364 3985 24392
rect 2372 24352 2378 24364
rect 3973 24361 3985 24364
rect 4019 24361 4031 24395
rect 3973 24355 4031 24361
rect 7006 24352 7012 24404
rect 7064 24392 7070 24404
rect 7101 24395 7159 24401
rect 7101 24392 7113 24395
rect 7064 24364 7113 24392
rect 7064 24352 7070 24364
rect 7101 24361 7113 24364
rect 7147 24361 7159 24395
rect 7926 24392 7932 24404
rect 7887 24364 7932 24392
rect 7101 24355 7159 24361
rect 7926 24352 7932 24364
rect 7984 24352 7990 24404
rect 10226 24352 10232 24404
rect 10284 24392 10290 24404
rect 10781 24395 10839 24401
rect 10781 24392 10793 24395
rect 10284 24364 10793 24392
rect 10284 24352 10290 24364
rect 10781 24361 10793 24364
rect 10827 24361 10839 24395
rect 10781 24355 10839 24361
rect 14182 24352 14188 24404
rect 14240 24392 14246 24404
rect 19702 24392 19708 24404
rect 14240 24364 15332 24392
rect 19663 24364 19708 24392
rect 14240 24352 14246 24364
rect 3418 24284 3424 24336
rect 3476 24324 3482 24336
rect 6273 24327 6331 24333
rect 6273 24324 6285 24327
rect 3476 24296 6285 24324
rect 3476 24284 3482 24296
rect 6273 24293 6285 24296
rect 6319 24293 6331 24327
rect 8754 24324 8760 24336
rect 6273 24287 6331 24293
rect 7208 24296 8760 24324
rect 1578 24256 1584 24268
rect 1539 24228 1584 24256
rect 1578 24216 1584 24228
rect 1636 24216 1642 24268
rect 4525 24259 4583 24265
rect 4525 24225 4537 24259
rect 4571 24256 4583 24259
rect 4890 24256 4896 24268
rect 4571 24228 4896 24256
rect 4571 24225 4583 24228
rect 4525 24219 4583 24225
rect 4890 24216 4896 24228
rect 4948 24216 4954 24268
rect 5994 24256 6000 24268
rect 5955 24228 6000 24256
rect 5994 24216 6000 24228
rect 6052 24216 6058 24268
rect 7006 24216 7012 24268
rect 7064 24256 7070 24268
rect 7208 24265 7236 24296
rect 8754 24284 8760 24296
rect 8812 24284 8818 24336
rect 15304 24324 15332 24364
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 20438 24392 20444 24404
rect 19935 24364 20444 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 20438 24352 20444 24364
rect 20496 24352 20502 24404
rect 20898 24392 20904 24404
rect 20859 24364 20904 24392
rect 20898 24352 20904 24364
rect 20956 24352 20962 24404
rect 21729 24395 21787 24401
rect 21008 24364 21680 24392
rect 19981 24327 20039 24333
rect 19981 24324 19993 24327
rect 15304 24296 19993 24324
rect 19981 24293 19993 24296
rect 20027 24324 20039 24327
rect 20070 24324 20076 24336
rect 20027 24296 20076 24324
rect 20027 24293 20039 24296
rect 19981 24287 20039 24293
rect 20070 24284 20076 24296
rect 20128 24324 20134 24336
rect 21008 24324 21036 24364
rect 20128 24296 21036 24324
rect 21085 24327 21143 24333
rect 20128 24284 20134 24296
rect 21085 24293 21097 24327
rect 21131 24293 21143 24327
rect 21085 24287 21143 24293
rect 7193 24259 7251 24265
rect 7193 24256 7205 24259
rect 7064 24228 7205 24256
rect 7064 24216 7070 24228
rect 7193 24225 7205 24228
rect 7239 24225 7251 24259
rect 7193 24219 7251 24225
rect 8018 24216 8024 24268
rect 8076 24256 8082 24268
rect 11333 24259 11391 24265
rect 11333 24256 11345 24259
rect 8076 24228 11345 24256
rect 8076 24216 8082 24228
rect 11333 24225 11345 24228
rect 11379 24225 11391 24259
rect 17589 24259 17647 24265
rect 11333 24219 11391 24225
rect 12406 24228 14412 24256
rect 1848 24191 1906 24197
rect 1848 24157 1860 24191
rect 1894 24188 1906 24191
rect 2222 24188 2228 24200
rect 1894 24160 2228 24188
rect 1894 24157 1906 24160
rect 1848 24151 1906 24157
rect 2222 24148 2228 24160
rect 2280 24148 2286 24200
rect 3142 24188 3148 24200
rect 2976 24160 3148 24188
rect 2976 24061 3004 24160
rect 3142 24148 3148 24160
rect 3200 24188 3206 24200
rect 4154 24191 4212 24197
rect 4154 24188 4166 24191
rect 3200 24160 4166 24188
rect 3200 24148 3206 24160
rect 4154 24157 4166 24160
rect 4200 24188 4212 24191
rect 4430 24188 4436 24200
rect 4200 24160 4436 24188
rect 4200 24157 4212 24160
rect 4154 24151 4212 24157
rect 4430 24148 4436 24160
rect 4488 24148 4494 24200
rect 4614 24148 4620 24200
rect 4672 24188 4678 24200
rect 6086 24188 6092 24200
rect 4672 24160 4717 24188
rect 6047 24160 6092 24188
rect 4672 24148 4678 24160
rect 6086 24148 6092 24160
rect 6144 24148 6150 24200
rect 7098 24188 7104 24200
rect 7059 24160 7104 24188
rect 7098 24148 7104 24160
rect 7156 24148 7162 24200
rect 8205 24191 8263 24197
rect 8205 24188 8217 24191
rect 7484 24160 8217 24188
rect 5629 24123 5687 24129
rect 5629 24089 5641 24123
rect 5675 24120 5687 24123
rect 5994 24120 6000 24132
rect 5675 24092 6000 24120
rect 5675 24089 5687 24092
rect 5629 24083 5687 24089
rect 5994 24080 6000 24092
rect 6052 24120 6058 24132
rect 6730 24120 6736 24132
rect 6052 24092 6736 24120
rect 6052 24080 6058 24092
rect 6730 24080 6736 24092
rect 6788 24080 6794 24132
rect 2961 24055 3019 24061
rect 2961 24021 2973 24055
rect 3007 24021 3019 24055
rect 2961 24015 3019 24021
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24052 4215 24055
rect 4522 24052 4528 24064
rect 4203 24024 4528 24052
rect 4203 24021 4215 24024
rect 4157 24015 4215 24021
rect 4522 24012 4528 24024
rect 4580 24052 4586 24064
rect 5350 24052 5356 24064
rect 4580 24024 5356 24052
rect 4580 24012 4586 24024
rect 5350 24012 5356 24024
rect 5408 24052 5414 24064
rect 7282 24052 7288 24064
rect 5408 24024 7288 24052
rect 5408 24012 5414 24024
rect 7282 24012 7288 24024
rect 7340 24012 7346 24064
rect 7484 24061 7512 24160
rect 8205 24157 8217 24160
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 9950 24148 9956 24200
rect 10008 24188 10014 24200
rect 10413 24191 10471 24197
rect 10413 24188 10425 24191
rect 10008 24160 10425 24188
rect 10008 24148 10014 24160
rect 10413 24157 10425 24160
rect 10459 24157 10471 24191
rect 12406 24188 12434 24228
rect 13446 24188 13452 24200
rect 10413 24151 10471 24157
rect 11440 24160 12434 24188
rect 13407 24160 13452 24188
rect 7929 24123 7987 24129
rect 7929 24089 7941 24123
rect 7975 24120 7987 24123
rect 8846 24120 8852 24132
rect 7975 24092 8852 24120
rect 7975 24089 7987 24092
rect 7929 24083 7987 24089
rect 8846 24080 8852 24092
rect 8904 24080 8910 24132
rect 10502 24080 10508 24132
rect 10560 24120 10566 24132
rect 10597 24123 10655 24129
rect 10597 24120 10609 24123
rect 10560 24092 10609 24120
rect 10560 24080 10566 24092
rect 10597 24089 10609 24092
rect 10643 24120 10655 24123
rect 11440 24120 11468 24160
rect 13446 24148 13452 24160
rect 13504 24148 13510 24200
rect 13725 24191 13783 24197
rect 13725 24157 13737 24191
rect 13771 24157 13783 24191
rect 13725 24151 13783 24157
rect 10643 24092 11468 24120
rect 11600 24123 11658 24129
rect 10643 24089 10655 24092
rect 10597 24083 10655 24089
rect 11600 24089 11612 24123
rect 11646 24120 11658 24123
rect 12158 24120 12164 24132
rect 11646 24092 12164 24120
rect 11646 24089 11658 24092
rect 11600 24083 11658 24089
rect 12158 24080 12164 24092
rect 12216 24080 12222 24132
rect 12986 24080 12992 24132
rect 13044 24120 13050 24132
rect 13633 24123 13691 24129
rect 13633 24120 13645 24123
rect 13044 24092 13645 24120
rect 13044 24080 13050 24092
rect 13633 24089 13645 24092
rect 13679 24089 13691 24123
rect 13633 24083 13691 24089
rect 7469 24055 7527 24061
rect 7469 24021 7481 24055
rect 7515 24021 7527 24055
rect 8110 24052 8116 24064
rect 8071 24024 8116 24052
rect 7469 24015 7527 24021
rect 8110 24012 8116 24024
rect 8168 24012 8174 24064
rect 8202 24012 8208 24064
rect 8260 24052 8266 24064
rect 12713 24055 12771 24061
rect 12713 24052 12725 24055
rect 8260 24024 12725 24052
rect 8260 24012 8266 24024
rect 12713 24021 12725 24024
rect 12759 24021 12771 24055
rect 13262 24052 13268 24064
rect 13223 24024 13268 24052
rect 12713 24015 12771 24021
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 13740 24052 13768 24151
rect 14090 24148 14096 24200
rect 14148 24188 14154 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 14148 24160 14289 24188
rect 14148 24148 14154 24160
rect 14277 24157 14289 24160
rect 14323 24157 14335 24191
rect 14384 24188 14412 24228
rect 17589 24225 17601 24259
rect 17635 24256 17647 24259
rect 19150 24256 19156 24268
rect 17635 24228 19156 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 14384 24160 16344 24188
rect 14277 24151 14335 24157
rect 14544 24123 14602 24129
rect 14544 24089 14556 24123
rect 14590 24120 14602 24123
rect 14918 24120 14924 24132
rect 14590 24092 14924 24120
rect 14590 24089 14602 24092
rect 14544 24083 14602 24089
rect 14918 24080 14924 24092
rect 14976 24080 14982 24132
rect 16316 24120 16344 24160
rect 16390 24148 16396 24200
rect 16448 24188 16454 24200
rect 16448 24160 16493 24188
rect 16448 24148 16454 24160
rect 16574 24148 16580 24200
rect 16632 24188 16638 24200
rect 16632 24160 16677 24188
rect 16632 24148 16638 24160
rect 17494 24148 17500 24200
rect 17552 24188 17558 24200
rect 17865 24191 17923 24197
rect 17865 24188 17877 24191
rect 17552 24160 17877 24188
rect 17552 24148 17558 24160
rect 17865 24157 17877 24160
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24188 19763 24191
rect 20346 24188 20352 24200
rect 19751 24160 20352 24188
rect 19751 24157 19763 24160
rect 19705 24151 19763 24157
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 20530 24188 20536 24200
rect 20491 24160 20536 24188
rect 20530 24148 20536 24160
rect 20588 24148 20594 24200
rect 21100 24188 21128 24287
rect 21652 24256 21680 24364
rect 21729 24361 21741 24395
rect 21775 24392 21787 24395
rect 22094 24392 22100 24404
rect 21775 24364 22100 24392
rect 21775 24361 21787 24364
rect 21729 24355 21787 24361
rect 22094 24352 22100 24364
rect 22152 24352 22158 24404
rect 22370 24352 22376 24404
rect 22428 24392 22434 24404
rect 23017 24395 23075 24401
rect 23017 24392 23029 24395
rect 22428 24364 23029 24392
rect 22428 24352 22434 24364
rect 23017 24361 23029 24364
rect 23063 24361 23075 24395
rect 23017 24355 23075 24361
rect 23750 24256 23756 24268
rect 21652 24228 23756 24256
rect 23750 24216 23756 24228
rect 23808 24256 23814 24268
rect 23845 24259 23903 24265
rect 23845 24256 23857 24259
rect 23808 24228 23857 24256
rect 23808 24216 23814 24228
rect 23845 24225 23857 24228
rect 23891 24225 23903 24259
rect 23845 24219 23903 24225
rect 21913 24191 21971 24197
rect 21913 24188 21925 24191
rect 21100 24160 21925 24188
rect 21913 24157 21925 24160
rect 21959 24157 21971 24191
rect 21913 24151 21971 24157
rect 23382 24148 23388 24200
rect 23440 24188 23446 24200
rect 23661 24191 23719 24197
rect 23661 24188 23673 24191
rect 23440 24160 23673 24188
rect 23440 24148 23446 24160
rect 23661 24157 23673 24160
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 19334 24120 19340 24132
rect 16316 24092 19340 24120
rect 19334 24080 19340 24092
rect 19392 24080 19398 24132
rect 20073 24123 20131 24129
rect 20073 24089 20085 24123
rect 20119 24120 20131 24123
rect 21266 24120 21272 24132
rect 20119 24092 21272 24120
rect 20119 24089 20131 24092
rect 20073 24083 20131 24089
rect 21266 24080 21272 24092
rect 21324 24080 21330 24132
rect 22925 24123 22983 24129
rect 22925 24089 22937 24123
rect 22971 24120 22983 24123
rect 23474 24120 23480 24132
rect 22971 24092 23480 24120
rect 22971 24089 22983 24092
rect 22925 24083 22983 24089
rect 23474 24080 23480 24092
rect 23532 24080 23538 24132
rect 15654 24052 15660 24064
rect 13740 24024 15660 24052
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 16298 24012 16304 24064
rect 16356 24052 16362 24064
rect 16485 24055 16543 24061
rect 16485 24052 16497 24055
rect 16356 24024 16497 24052
rect 16356 24012 16362 24024
rect 16485 24021 16497 24024
rect 16531 24021 16543 24055
rect 16485 24015 16543 24021
rect 16758 24012 16764 24064
rect 16816 24052 16822 24064
rect 20901 24055 20959 24061
rect 20901 24052 20913 24055
rect 16816 24024 20913 24052
rect 16816 24012 16822 24024
rect 20901 24021 20913 24024
rect 20947 24021 20959 24055
rect 20901 24015 20959 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 3234 23808 3240 23860
rect 3292 23848 3298 23860
rect 3694 23848 3700 23860
rect 3292 23820 3700 23848
rect 3292 23808 3298 23820
rect 3694 23808 3700 23820
rect 3752 23848 3758 23860
rect 4617 23851 4675 23857
rect 4617 23848 4629 23851
rect 3752 23820 4629 23848
rect 3752 23808 3758 23820
rect 4617 23817 4629 23820
rect 4663 23817 4675 23851
rect 5994 23848 6000 23860
rect 5955 23820 6000 23848
rect 4617 23811 4675 23817
rect 5994 23808 6000 23820
rect 6052 23808 6058 23860
rect 6086 23808 6092 23860
rect 6144 23848 6150 23860
rect 6917 23851 6975 23857
rect 6917 23848 6929 23851
rect 6144 23820 6929 23848
rect 6144 23808 6150 23820
rect 6917 23817 6929 23820
rect 6963 23817 6975 23851
rect 6917 23811 6975 23817
rect 7929 23851 7987 23857
rect 7929 23817 7941 23851
rect 7975 23848 7987 23851
rect 8110 23848 8116 23860
rect 7975 23820 8116 23848
rect 7975 23817 7987 23820
rect 7929 23811 7987 23817
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 9766 23848 9772 23860
rect 9727 23820 9772 23848
rect 9766 23808 9772 23820
rect 9824 23808 9830 23860
rect 12158 23848 12164 23860
rect 12119 23820 12164 23848
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 14182 23848 14188 23860
rect 12268 23820 14188 23848
rect 3602 23780 3608 23792
rect 2516 23752 3608 23780
rect 2516 23721 2544 23752
rect 3602 23740 3608 23752
rect 3660 23740 3666 23792
rect 5169 23783 5227 23789
rect 5169 23749 5181 23783
rect 5215 23780 5227 23783
rect 6733 23783 6791 23789
rect 6733 23780 6745 23783
rect 5215 23752 6745 23780
rect 5215 23749 5227 23752
rect 5169 23743 5227 23749
rect 2501 23715 2559 23721
rect 2501 23681 2513 23715
rect 2547 23681 2559 23715
rect 2501 23675 2559 23681
rect 2685 23715 2743 23721
rect 2685 23681 2697 23715
rect 2731 23712 2743 23715
rect 3234 23712 3240 23724
rect 2731 23684 3240 23712
rect 2731 23681 2743 23684
rect 2685 23675 2743 23681
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 3329 23715 3387 23721
rect 3329 23681 3341 23715
rect 3375 23681 3387 23715
rect 3329 23675 3387 23681
rect 4157 23715 4215 23721
rect 4157 23681 4169 23715
rect 4203 23712 4215 23715
rect 4706 23712 4712 23724
rect 4203 23684 4712 23712
rect 4203 23681 4215 23684
rect 4157 23675 4215 23681
rect 2593 23647 2651 23653
rect 2593 23613 2605 23647
rect 2639 23644 2651 23647
rect 3344 23644 3372 23675
rect 4706 23672 4712 23684
rect 4764 23712 4770 23724
rect 6012 23721 6040 23752
rect 6733 23749 6745 23752
rect 6779 23780 6791 23783
rect 8202 23780 8208 23792
rect 6779 23752 8208 23780
rect 6779 23749 6791 23752
rect 6733 23743 6791 23749
rect 8202 23740 8208 23752
rect 8260 23740 8266 23792
rect 9674 23780 9680 23792
rect 8588 23752 9680 23780
rect 5353 23715 5411 23721
rect 5353 23712 5365 23715
rect 4764 23684 5365 23712
rect 4764 23672 4770 23684
rect 5353 23681 5365 23684
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23681 5871 23715
rect 5813 23675 5871 23681
rect 5997 23715 6055 23721
rect 5997 23681 6009 23715
rect 6043 23681 6055 23715
rect 5997 23675 6055 23681
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 2639 23616 3372 23644
rect 2639 23613 2651 23616
rect 2593 23607 2651 23613
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 3697 23647 3755 23653
rect 3476 23616 3521 23644
rect 3476 23604 3482 23616
rect 3697 23613 3709 23647
rect 3743 23644 3755 23647
rect 4614 23644 4620 23656
rect 3743 23616 4620 23644
rect 3743 23613 3755 23616
rect 3697 23607 3755 23613
rect 4614 23604 4620 23616
rect 4672 23604 4678 23656
rect 5828 23644 5856 23675
rect 6564 23644 6592 23675
rect 7282 23672 7288 23724
rect 7340 23712 7346 23724
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 7340 23684 7757 23712
rect 7340 23672 7346 23684
rect 7745 23681 7757 23684
rect 7791 23681 7803 23715
rect 7745 23675 7803 23681
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23712 7987 23715
rect 8588 23712 8616 23752
rect 9674 23740 9680 23752
rect 9732 23740 9738 23792
rect 12268 23780 12296 23820
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 14274 23808 14280 23860
rect 14332 23848 14338 23860
rect 14461 23851 14519 23857
rect 14332 23820 14377 23848
rect 14332 23808 14338 23820
rect 14461 23817 14473 23851
rect 14507 23817 14519 23851
rect 14918 23848 14924 23860
rect 14879 23820 14924 23848
rect 14461 23811 14519 23817
rect 13265 23783 13323 23789
rect 13265 23780 13277 23783
rect 10796 23752 12296 23780
rect 12360 23752 13277 23780
rect 8662 23721 8668 23724
rect 7975 23684 8616 23712
rect 7975 23681 7987 23684
rect 7929 23675 7987 23681
rect 8656 23675 8668 23721
rect 8720 23712 8726 23724
rect 10796 23721 10824 23752
rect 12360 23721 12388 23752
rect 13265 23749 13277 23752
rect 13311 23749 13323 23783
rect 13265 23743 13323 23749
rect 10781 23715 10839 23721
rect 8720 23684 8756 23712
rect 7944 23644 7972 23675
rect 8662 23672 8668 23675
rect 8720 23672 8726 23684
rect 10781 23681 10793 23715
rect 10827 23681 10839 23715
rect 10781 23675 10839 23681
rect 12345 23715 12403 23721
rect 12345 23681 12357 23715
rect 12391 23681 12403 23715
rect 12345 23675 12403 23681
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23712 12495 23715
rect 12526 23712 12532 23724
rect 12483 23684 12532 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 12526 23672 12532 23684
rect 12584 23672 12590 23724
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 12713 23715 12771 23721
rect 12713 23681 12725 23715
rect 12759 23712 12771 23715
rect 12802 23712 12808 23724
rect 12759 23684 12808 23712
rect 12759 23681 12771 23684
rect 12713 23675 12771 23681
rect 5828 23616 7972 23644
rect 8018 23604 8024 23656
rect 8076 23644 8082 23656
rect 8389 23647 8447 23653
rect 8389 23644 8401 23647
rect 8076 23616 8401 23644
rect 8076 23604 8082 23616
rect 8389 23613 8401 23616
rect 8435 23613 8447 23647
rect 8389 23607 8447 23613
rect 10689 23647 10747 23653
rect 10689 23613 10701 23647
rect 10735 23613 10747 23647
rect 12636 23644 12664 23675
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 13170 23712 13176 23724
rect 13131 23684 13176 23712
rect 13170 23672 13176 23684
rect 13228 23672 13234 23724
rect 13354 23712 13360 23724
rect 13315 23684 13360 23712
rect 13354 23672 13360 23684
rect 13412 23672 13418 23724
rect 14476 23712 14504 23811
rect 14918 23808 14924 23820
rect 14976 23808 14982 23860
rect 16206 23848 16212 23860
rect 16119 23820 16212 23848
rect 16206 23808 16212 23820
rect 16264 23848 16270 23860
rect 16482 23848 16488 23860
rect 16264 23820 16488 23848
rect 16264 23808 16270 23820
rect 16482 23808 16488 23820
rect 16540 23808 16546 23860
rect 18230 23848 18236 23860
rect 18191 23820 18236 23848
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 20714 23808 20720 23860
rect 20772 23848 20778 23860
rect 22205 23851 22263 23857
rect 22205 23848 22217 23851
rect 20772 23820 22217 23848
rect 20772 23808 20778 23820
rect 22205 23817 22217 23820
rect 22251 23817 22263 23851
rect 22205 23811 22263 23817
rect 23293 23851 23351 23857
rect 23293 23817 23305 23851
rect 23339 23848 23351 23851
rect 23382 23848 23388 23860
rect 23339 23820 23388 23848
rect 23339 23817 23351 23820
rect 23293 23811 23351 23817
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 20990 23780 20996 23792
rect 16500 23752 20996 23780
rect 15105 23715 15163 23721
rect 15105 23712 15117 23715
rect 14476 23684 15117 23712
rect 15105 23681 15117 23684
rect 15151 23681 15163 23715
rect 16022 23712 16028 23724
rect 15983 23684 16028 23712
rect 15105 23675 15163 23681
rect 16022 23672 16028 23684
rect 16080 23672 16086 23724
rect 16298 23712 16304 23724
rect 16259 23684 16304 23712
rect 16298 23672 16304 23684
rect 16356 23672 16362 23724
rect 13446 23644 13452 23656
rect 12636 23616 13452 23644
rect 10689 23607 10747 23613
rect 4430 23508 4436 23520
rect 4343 23480 4436 23508
rect 4430 23468 4436 23480
rect 4488 23508 4494 23520
rect 4798 23508 4804 23520
rect 4488 23480 4804 23508
rect 4488 23468 4494 23480
rect 4798 23468 4804 23480
rect 4856 23508 4862 23520
rect 10704 23508 10732 23607
rect 13446 23604 13452 23616
rect 13504 23604 13510 23656
rect 16500 23644 16528 23752
rect 20990 23740 20996 23752
rect 21048 23740 21054 23792
rect 22002 23780 22008 23792
rect 21963 23752 22008 23780
rect 22002 23740 22008 23752
rect 22060 23740 22066 23792
rect 17109 23715 17167 23721
rect 17109 23712 17121 23715
rect 13740 23616 16528 23644
rect 16592 23684 17121 23712
rect 11882 23536 11888 23588
rect 11940 23576 11946 23588
rect 13740 23576 13768 23616
rect 13906 23576 13912 23588
rect 11940 23548 13768 23576
rect 13867 23548 13912 23576
rect 11940 23536 11946 23548
rect 13906 23536 13912 23548
rect 13964 23536 13970 23588
rect 14090 23536 14096 23588
rect 14148 23576 14154 23588
rect 16025 23579 16083 23585
rect 14148 23548 15976 23576
rect 14148 23536 14154 23548
rect 11146 23508 11152 23520
rect 4856 23480 10732 23508
rect 11107 23480 11152 23508
rect 4856 23468 4862 23480
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 13262 23468 13268 23520
rect 13320 23508 13326 23520
rect 14277 23511 14335 23517
rect 14277 23508 14289 23511
rect 13320 23480 14289 23508
rect 13320 23468 13326 23480
rect 14277 23477 14289 23480
rect 14323 23477 14335 23511
rect 15948 23508 15976 23548
rect 16025 23545 16037 23579
rect 16071 23576 16083 23579
rect 16592 23576 16620 23684
rect 17109 23681 17121 23684
rect 17155 23681 17167 23715
rect 17109 23675 17167 23681
rect 20530 23672 20536 23724
rect 20588 23712 20594 23724
rect 23198 23712 23204 23724
rect 20588 23684 21404 23712
rect 23159 23684 23204 23712
rect 20588 23672 20594 23684
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 16071 23548 16620 23576
rect 16684 23616 16865 23644
rect 16071 23545 16083 23548
rect 16025 23539 16083 23545
rect 16684 23508 16712 23616
rect 16853 23613 16865 23616
rect 16899 23613 16911 23647
rect 18690 23644 18696 23656
rect 18651 23616 18696 23644
rect 16853 23607 16911 23613
rect 18690 23604 18696 23616
rect 18748 23604 18754 23656
rect 18969 23647 19027 23653
rect 18969 23613 18981 23647
rect 19015 23644 19027 23647
rect 19150 23644 19156 23656
rect 19015 23616 19156 23644
rect 19015 23613 19027 23616
rect 18969 23607 19027 23613
rect 19150 23604 19156 23616
rect 19208 23604 19214 23656
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 20625 23647 20683 23653
rect 20625 23644 20637 23647
rect 19392 23616 20637 23644
rect 19392 23604 19398 23616
rect 20625 23613 20637 23616
rect 20671 23613 20683 23647
rect 20625 23607 20683 23613
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23644 20959 23647
rect 21266 23644 21272 23656
rect 20947 23616 21272 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 20640 23576 20668 23607
rect 21266 23604 21272 23616
rect 21324 23604 21330 23656
rect 21376 23644 21404 23684
rect 23198 23672 23204 23684
rect 23256 23672 23262 23724
rect 23290 23672 23296 23724
rect 23348 23712 23354 23724
rect 23385 23715 23443 23721
rect 23385 23712 23397 23715
rect 23348 23684 23397 23712
rect 23348 23672 23354 23684
rect 23385 23681 23397 23684
rect 23431 23712 23443 23715
rect 23934 23712 23940 23724
rect 23431 23684 23940 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 23934 23672 23940 23684
rect 23992 23672 23998 23724
rect 23569 23647 23627 23653
rect 23569 23644 23581 23647
rect 21376 23616 23581 23644
rect 23569 23613 23581 23616
rect 23615 23613 23627 23647
rect 23569 23607 23627 23613
rect 22462 23576 22468 23588
rect 20640 23548 22468 23576
rect 22462 23536 22468 23548
rect 22520 23536 22526 23588
rect 23017 23579 23075 23585
rect 23017 23545 23029 23579
rect 23063 23576 23075 23579
rect 23474 23576 23480 23588
rect 23063 23548 23480 23576
rect 23063 23545 23075 23548
rect 23017 23539 23075 23545
rect 23474 23536 23480 23548
rect 23532 23536 23538 23588
rect 15948 23480 16712 23508
rect 14277 23471 14335 23477
rect 20990 23468 20996 23520
rect 21048 23508 21054 23520
rect 22189 23511 22247 23517
rect 22189 23508 22201 23511
rect 21048 23480 22201 23508
rect 21048 23468 21054 23480
rect 22189 23477 22201 23480
rect 22235 23477 22247 23511
rect 22370 23508 22376 23520
rect 22331 23480 22376 23508
rect 22189 23471 22247 23477
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 8573 23307 8631 23313
rect 8573 23273 8585 23307
rect 8619 23304 8631 23307
rect 8662 23304 8668 23316
rect 8619 23276 8668 23304
rect 8619 23273 8631 23276
rect 8573 23267 8631 23273
rect 8662 23264 8668 23276
rect 8720 23264 8726 23316
rect 8846 23264 8852 23316
rect 8904 23304 8910 23316
rect 12802 23304 12808 23316
rect 8904 23276 12808 23304
rect 8904 23264 8910 23276
rect 12802 23264 12808 23276
rect 12860 23304 12866 23316
rect 12989 23307 13047 23313
rect 12989 23304 13001 23307
rect 12860 23276 13001 23304
rect 12860 23264 12866 23276
rect 12989 23273 13001 23276
rect 13035 23273 13047 23307
rect 12989 23267 13047 23273
rect 16022 23264 16028 23316
rect 16080 23304 16086 23316
rect 16301 23307 16359 23313
rect 16301 23304 16313 23307
rect 16080 23276 16313 23304
rect 16080 23264 16086 23276
rect 16301 23273 16313 23276
rect 16347 23273 16359 23307
rect 16301 23267 16359 23273
rect 18138 23264 18144 23316
rect 18196 23304 18202 23316
rect 18598 23304 18604 23316
rect 18196 23276 18604 23304
rect 18196 23264 18202 23276
rect 18598 23264 18604 23276
rect 18656 23304 18662 23316
rect 18877 23307 18935 23313
rect 18877 23304 18889 23307
rect 18656 23276 18889 23304
rect 18656 23264 18662 23276
rect 18877 23273 18889 23276
rect 18923 23273 18935 23307
rect 18877 23267 18935 23273
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 19981 23307 20039 23313
rect 19981 23304 19993 23307
rect 19484 23276 19993 23304
rect 19484 23264 19490 23276
rect 19981 23273 19993 23276
rect 20027 23273 20039 23307
rect 20898 23304 20904 23316
rect 20859 23276 20904 23304
rect 19981 23267 20039 23273
rect 20898 23264 20904 23276
rect 20956 23264 20962 23316
rect 23934 23304 23940 23316
rect 23895 23276 23940 23304
rect 23934 23264 23940 23276
rect 23992 23264 23998 23316
rect 4249 23239 4307 23245
rect 4249 23205 4261 23239
rect 4295 23236 4307 23239
rect 4798 23236 4804 23248
rect 4295 23208 4804 23236
rect 4295 23205 4307 23208
rect 4249 23199 4307 23205
rect 4798 23196 4804 23208
rect 4856 23196 4862 23248
rect 6546 23236 6552 23248
rect 6507 23208 6552 23236
rect 6546 23196 6552 23208
rect 6604 23196 6610 23248
rect 8389 23239 8447 23245
rect 8389 23205 8401 23239
rect 8435 23236 8447 23239
rect 9309 23239 9367 23245
rect 9309 23236 9321 23239
rect 8435 23208 9321 23236
rect 8435 23205 8447 23208
rect 8389 23199 8447 23205
rect 9309 23205 9321 23208
rect 9355 23205 9367 23239
rect 9309 23199 9367 23205
rect 3973 23171 4031 23177
rect 3973 23137 3985 23171
rect 4019 23168 4031 23171
rect 4338 23168 4344 23180
rect 4019 23140 4344 23168
rect 4019 23137 4031 23140
rect 3973 23131 4031 23137
rect 4338 23128 4344 23140
rect 4396 23168 4402 23180
rect 4706 23168 4712 23180
rect 4396 23140 4712 23168
rect 4396 23128 4402 23140
rect 4706 23128 4712 23140
rect 4764 23128 4770 23180
rect 5166 23168 5172 23180
rect 5000 23140 5172 23168
rect 5000 23109 5028 23140
rect 5166 23128 5172 23140
rect 5224 23168 5230 23180
rect 15378 23168 15384 23180
rect 5224 23140 12434 23168
rect 15339 23140 15384 23168
rect 5224 23128 5230 23140
rect 4985 23103 5043 23109
rect 4985 23069 4997 23103
rect 5031 23069 5043 23103
rect 4985 23063 5043 23069
rect 5350 23060 5356 23112
rect 5408 23100 5414 23112
rect 5905 23103 5963 23109
rect 5905 23100 5917 23103
rect 5408 23072 5917 23100
rect 5408 23060 5414 23072
rect 5905 23069 5917 23072
rect 5951 23069 5963 23103
rect 6086 23100 6092 23112
rect 6047 23072 6092 23100
rect 5905 23063 5963 23069
rect 6086 23060 6092 23072
rect 6144 23060 6150 23112
rect 6825 23103 6883 23109
rect 6825 23069 6837 23103
rect 6871 23100 6883 23103
rect 7098 23100 7104 23112
rect 6871 23072 7104 23100
rect 6871 23069 6883 23072
rect 6825 23063 6883 23069
rect 7098 23060 7104 23072
rect 7156 23060 7162 23112
rect 8481 23103 8539 23109
rect 8481 23100 8493 23103
rect 8036 23072 8493 23100
rect 6549 23035 6607 23041
rect 6549 23001 6561 23035
rect 6595 23032 6607 23035
rect 8036 23032 8064 23072
rect 8481 23069 8493 23072
rect 8527 23100 8539 23103
rect 8846 23100 8852 23112
rect 8527 23072 8852 23100
rect 8527 23069 8539 23072
rect 8481 23063 8539 23069
rect 8846 23060 8852 23072
rect 8904 23060 8910 23112
rect 9582 23100 9588 23112
rect 9543 23072 9588 23100
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 6595 23004 8064 23032
rect 8113 23035 8171 23041
rect 6595 23001 6607 23004
rect 6549 22995 6607 23001
rect 8113 23001 8125 23035
rect 8159 23032 8171 23035
rect 8386 23032 8392 23044
rect 8159 23004 8392 23032
rect 8159 23001 8171 23004
rect 8113 22995 8171 23001
rect 8386 22992 8392 23004
rect 8444 22992 8450 23044
rect 9309 23035 9367 23041
rect 9309 23001 9321 23035
rect 9355 23032 9367 23035
rect 10226 23032 10232 23044
rect 9355 23004 10232 23032
rect 9355 23001 9367 23004
rect 9309 22995 9367 23001
rect 10226 22992 10232 23004
rect 10284 22992 10290 23044
rect 12406 23032 12434 23140
rect 15378 23128 15384 23140
rect 15436 23128 15442 23180
rect 15841 23171 15899 23177
rect 15841 23137 15853 23171
rect 15887 23168 15899 23171
rect 15930 23168 15936 23180
rect 15887 23140 15936 23168
rect 15887 23137 15899 23140
rect 15841 23131 15899 23137
rect 15930 23128 15936 23140
rect 15988 23128 15994 23180
rect 16574 23168 16580 23180
rect 16487 23140 16580 23168
rect 16574 23128 16580 23140
rect 16632 23168 16638 23180
rect 17402 23168 17408 23180
rect 16632 23140 17408 23168
rect 16632 23128 16638 23140
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 19392 23140 19441 23168
rect 19392 23128 19398 23140
rect 19429 23137 19441 23140
rect 19475 23137 19487 23171
rect 19429 23131 19487 23137
rect 20438 23128 20444 23180
rect 20496 23168 20502 23180
rect 20898 23168 20904 23180
rect 20496 23140 20904 23168
rect 20496 23128 20502 23140
rect 20898 23128 20904 23140
rect 20956 23168 20962 23180
rect 21085 23171 21143 23177
rect 21085 23168 21097 23171
rect 20956 23140 21097 23168
rect 20956 23128 20962 23140
rect 21085 23137 21097 23140
rect 21131 23137 21143 23171
rect 21085 23131 21143 23137
rect 21177 23171 21235 23177
rect 21177 23137 21189 23171
rect 21223 23168 21235 23171
rect 21726 23168 21732 23180
rect 21223 23140 21732 23168
rect 21223 23137 21235 23140
rect 21177 23131 21235 23137
rect 21726 23128 21732 23140
rect 21784 23128 21790 23180
rect 22186 23128 22192 23180
rect 22244 23168 22250 23180
rect 22557 23171 22615 23177
rect 22557 23168 22569 23171
rect 22244 23140 22569 23168
rect 22244 23128 22250 23140
rect 22557 23137 22569 23140
rect 22603 23137 22615 23171
rect 22557 23131 22615 23137
rect 15102 23060 15108 23112
rect 15160 23100 15166 23112
rect 15473 23103 15531 23109
rect 15473 23100 15485 23103
rect 15160 23072 15485 23100
rect 15160 23060 15166 23072
rect 15473 23069 15485 23072
rect 15519 23069 15531 23103
rect 15473 23063 15531 23069
rect 16390 23060 16396 23112
rect 16448 23100 16454 23112
rect 16485 23103 16543 23109
rect 16485 23100 16497 23103
rect 16448 23072 16497 23100
rect 16448 23060 16454 23072
rect 16485 23069 16497 23072
rect 16531 23069 16543 23103
rect 16485 23063 16543 23069
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 12897 23035 12955 23041
rect 12897 23032 12909 23035
rect 12406 23004 12909 23032
rect 12897 23001 12909 23004
rect 12943 23032 12955 23035
rect 16574 23032 16580 23044
rect 12943 23004 16580 23032
rect 12943 23001 12955 23004
rect 12897 22995 12955 23001
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 16684 23032 16712 23063
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17494 23100 17500 23112
rect 16816 23072 16861 23100
rect 17455 23072 17500 23100
rect 16816 23060 16822 23072
rect 17494 23060 17500 23072
rect 17552 23060 17558 23112
rect 19797 23103 19855 23109
rect 19797 23100 19809 23103
rect 19444 23072 19809 23100
rect 19444 23044 19472 23072
rect 19797 23069 19809 23072
rect 19843 23069 19855 23103
rect 19797 23063 19855 23069
rect 16684 23004 16979 23032
rect 3418 22924 3424 22976
rect 3476 22964 3482 22976
rect 4433 22967 4491 22973
rect 4433 22964 4445 22967
rect 3476 22936 4445 22964
rect 3476 22924 3482 22936
rect 4433 22933 4445 22936
rect 4479 22933 4491 22967
rect 4433 22927 4491 22933
rect 4890 22924 4896 22976
rect 4948 22964 4954 22976
rect 5077 22967 5135 22973
rect 5077 22964 5089 22967
rect 4948 22936 5089 22964
rect 4948 22924 4954 22936
rect 5077 22933 5089 22936
rect 5123 22933 5135 22967
rect 5077 22927 5135 22933
rect 6089 22967 6147 22973
rect 6089 22933 6101 22967
rect 6135 22964 6147 22967
rect 6733 22967 6791 22973
rect 6733 22964 6745 22967
rect 6135 22936 6745 22964
rect 6135 22933 6147 22936
rect 6089 22927 6147 22933
rect 6733 22933 6745 22936
rect 6779 22933 6791 22967
rect 6733 22927 6791 22933
rect 7834 22924 7840 22976
rect 7892 22964 7898 22976
rect 8205 22967 8263 22973
rect 8205 22964 8217 22967
rect 7892 22936 8217 22964
rect 7892 22924 7898 22936
rect 8205 22933 8217 22936
rect 8251 22933 8263 22967
rect 8205 22927 8263 22933
rect 9398 22924 9404 22976
rect 9456 22964 9462 22976
rect 9493 22967 9551 22973
rect 9493 22964 9505 22967
rect 9456 22936 9505 22964
rect 9456 22924 9462 22936
rect 9493 22933 9505 22936
rect 9539 22933 9551 22967
rect 9493 22927 9551 22933
rect 14458 22924 14464 22976
rect 14516 22964 14522 22976
rect 15102 22964 15108 22976
rect 14516 22936 15108 22964
rect 14516 22924 14522 22936
rect 15102 22924 15108 22936
rect 15160 22924 15166 22976
rect 15838 22924 15844 22976
rect 15896 22964 15902 22976
rect 16114 22964 16120 22976
rect 15896 22936 16120 22964
rect 15896 22924 15902 22936
rect 16114 22924 16120 22936
rect 16172 22924 16178 22976
rect 16951 22964 16979 23004
rect 17126 22992 17132 23044
rect 17184 23032 17190 23044
rect 17742 23035 17800 23041
rect 17742 23032 17754 23035
rect 17184 23004 17754 23032
rect 17184 22992 17190 23004
rect 17742 23001 17754 23004
rect 17788 23001 17800 23035
rect 17742 22995 17800 23001
rect 19426 22992 19432 23044
rect 19484 22992 19490 23044
rect 19705 23035 19763 23041
rect 19705 23001 19717 23035
rect 19751 23032 19763 23035
rect 20254 23032 20260 23044
rect 19751 23004 20260 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 20254 22992 20260 23004
rect 20312 23032 20318 23044
rect 20456 23032 20484 23128
rect 21266 23100 21272 23112
rect 21227 23072 21272 23100
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 21361 23103 21419 23109
rect 21361 23069 21373 23103
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 22097 23103 22155 23109
rect 22097 23069 22109 23103
rect 22143 23100 22155 23103
rect 22370 23100 22376 23112
rect 22143 23072 22376 23100
rect 22143 23069 22155 23072
rect 22097 23063 22155 23069
rect 20312 23004 20484 23032
rect 20312 22992 20318 23004
rect 17954 22964 17960 22976
rect 16951 22936 17960 22964
rect 17954 22924 17960 22936
rect 18012 22924 18018 22976
rect 19613 22967 19671 22973
rect 19613 22933 19625 22967
rect 19659 22964 19671 22967
rect 20070 22964 20076 22976
rect 19659 22936 20076 22964
rect 19659 22933 19671 22936
rect 19613 22927 19671 22933
rect 20070 22924 20076 22936
rect 20128 22964 20134 22976
rect 21376 22964 21404 23063
rect 22370 23060 22376 23072
rect 22428 23060 22434 23112
rect 22802 23035 22860 23041
rect 22802 23032 22814 23035
rect 22066 23004 22814 23032
rect 20128 22936 21404 22964
rect 21913 22967 21971 22973
rect 20128 22924 20134 22936
rect 21913 22933 21925 22967
rect 21959 22964 21971 22967
rect 22066 22964 22094 23004
rect 22802 23001 22814 23004
rect 22848 23001 22860 23035
rect 22802 22995 22860 23001
rect 21959 22936 22094 22964
rect 21959 22933 21971 22936
rect 21913 22927 21971 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22760 3663 22763
rect 3694 22760 3700 22772
rect 3651 22732 3700 22760
rect 3651 22729 3663 22732
rect 3605 22723 3663 22729
rect 3694 22720 3700 22732
rect 3752 22720 3758 22772
rect 5537 22763 5595 22769
rect 5537 22729 5549 22763
rect 5583 22760 5595 22763
rect 5902 22760 5908 22772
rect 5583 22732 5908 22760
rect 5583 22729 5595 22732
rect 5537 22723 5595 22729
rect 5902 22720 5908 22732
rect 5960 22720 5966 22772
rect 10226 22760 10232 22772
rect 10187 22732 10232 22760
rect 10226 22720 10232 22732
rect 10284 22720 10290 22772
rect 15562 22760 15568 22772
rect 15523 22732 15568 22760
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 16758 22760 16764 22772
rect 16632 22732 16764 22760
rect 16632 22720 16638 22732
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 17126 22760 17132 22772
rect 17087 22732 17132 22760
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17402 22720 17408 22772
rect 17460 22760 17466 22772
rect 18785 22763 18843 22769
rect 18785 22760 18797 22763
rect 17460 22732 18797 22760
rect 17460 22720 17466 22732
rect 18785 22729 18797 22732
rect 18831 22760 18843 22763
rect 18966 22760 18972 22772
rect 18831 22732 18972 22760
rect 18831 22729 18843 22732
rect 18785 22723 18843 22729
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 20073 22763 20131 22769
rect 20073 22729 20085 22763
rect 20119 22760 20131 22763
rect 20714 22760 20720 22772
rect 20119 22732 20720 22760
rect 20119 22729 20131 22732
rect 20073 22723 20131 22729
rect 20714 22720 20720 22732
rect 20772 22720 20778 22772
rect 23474 22720 23480 22772
rect 23532 22760 23538 22772
rect 23569 22763 23627 22769
rect 23569 22760 23581 22763
rect 23532 22732 23581 22760
rect 23532 22720 23538 22732
rect 23569 22729 23581 22732
rect 23615 22729 23627 22763
rect 23569 22723 23627 22729
rect 3418 22692 3424 22704
rect 3379 22664 3424 22692
rect 3418 22652 3424 22664
rect 3476 22652 3482 22704
rect 5810 22692 5816 22704
rect 5368 22664 5816 22692
rect 2774 22584 2780 22636
rect 2832 22624 2838 22636
rect 2958 22624 2964 22636
rect 2832 22596 2877 22624
rect 2919 22596 2964 22624
rect 2832 22584 2838 22596
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 3697 22627 3755 22633
rect 3697 22624 3709 22627
rect 3568 22596 3709 22624
rect 3568 22584 3574 22596
rect 3697 22593 3709 22596
rect 3743 22593 3755 22627
rect 3697 22587 3755 22593
rect 4157 22627 4215 22633
rect 4157 22593 4169 22627
rect 4203 22593 4215 22627
rect 4338 22624 4344 22636
rect 4299 22596 4344 22624
rect 4157 22587 4215 22593
rect 4172 22556 4200 22587
rect 4338 22584 4344 22596
rect 4396 22624 4402 22636
rect 4614 22624 4620 22636
rect 4396 22596 4620 22624
rect 4396 22584 4402 22596
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 4798 22584 4804 22636
rect 4856 22624 4862 22636
rect 5368 22633 5396 22664
rect 5810 22652 5816 22664
rect 5868 22652 5874 22704
rect 6546 22652 6552 22704
rect 6604 22692 6610 22704
rect 6794 22695 6852 22701
rect 6794 22692 6806 22695
rect 6604 22664 6806 22692
rect 6604 22652 6610 22664
rect 6794 22661 6806 22664
rect 6840 22661 6852 22695
rect 11146 22692 11152 22704
rect 6794 22655 6852 22661
rect 10520 22664 11152 22692
rect 5353 22627 5411 22633
rect 5353 22624 5365 22627
rect 4856 22596 5365 22624
rect 4856 22584 4862 22596
rect 5353 22593 5365 22596
rect 5399 22593 5411 22627
rect 5353 22587 5411 22593
rect 5537 22627 5595 22633
rect 5537 22593 5549 22627
rect 5583 22624 5595 22627
rect 6454 22624 6460 22636
rect 5583 22596 6460 22624
rect 5583 22593 5595 22596
rect 5537 22587 5595 22593
rect 6454 22584 6460 22596
rect 6512 22584 6518 22636
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22624 9459 22627
rect 9490 22624 9496 22636
rect 9447 22596 9496 22624
rect 9447 22593 9459 22596
rect 9401 22587 9459 22593
rect 9490 22584 9496 22596
rect 9548 22584 9554 22636
rect 10520 22633 10548 22664
rect 11146 22652 11152 22664
rect 11204 22692 11210 22704
rect 11793 22695 11851 22701
rect 11793 22692 11805 22695
rect 11204 22664 11805 22692
rect 11204 22652 11210 22664
rect 11793 22661 11805 22664
rect 11839 22661 11851 22695
rect 11793 22655 11851 22661
rect 12250 22652 12256 22704
rect 12308 22692 12314 22704
rect 15473 22695 15531 22701
rect 12308 22664 12434 22692
rect 12308 22652 12314 22664
rect 10413 22627 10471 22633
rect 10413 22624 10425 22627
rect 9784 22596 10425 22624
rect 4982 22556 4988 22568
rect 4172 22528 4988 22556
rect 4982 22516 4988 22528
rect 5040 22516 5046 22568
rect 5442 22516 5448 22568
rect 5500 22556 5506 22568
rect 6549 22559 6607 22565
rect 6549 22556 6561 22559
rect 5500 22528 6561 22556
rect 5500 22516 5506 22528
rect 6549 22525 6561 22528
rect 6595 22525 6607 22559
rect 6549 22519 6607 22525
rect 9309 22559 9367 22565
rect 9309 22525 9321 22559
rect 9355 22556 9367 22559
rect 9355 22528 9444 22556
rect 9355 22525 9367 22528
rect 9309 22519 9367 22525
rect 2682 22448 2688 22500
rect 2740 22488 2746 22500
rect 4154 22488 4160 22500
rect 2740 22460 4016 22488
rect 4115 22460 4160 22488
rect 2740 22448 2746 22460
rect 2866 22420 2872 22432
rect 2827 22392 2872 22420
rect 2866 22380 2872 22392
rect 2924 22380 2930 22432
rect 3326 22380 3332 22432
rect 3384 22420 3390 22432
rect 3421 22423 3479 22429
rect 3421 22420 3433 22423
rect 3384 22392 3433 22420
rect 3384 22380 3390 22392
rect 3421 22389 3433 22392
rect 3467 22389 3479 22423
rect 3988 22420 4016 22460
rect 4154 22448 4160 22460
rect 4212 22448 4218 22500
rect 4338 22420 4344 22432
rect 3988 22392 4344 22420
rect 3421 22383 3479 22389
rect 4338 22380 4344 22392
rect 4396 22380 4402 22432
rect 7834 22380 7840 22432
rect 7892 22420 7898 22432
rect 7929 22423 7987 22429
rect 7929 22420 7941 22423
rect 7892 22392 7941 22420
rect 7892 22380 7898 22392
rect 7929 22389 7941 22392
rect 7975 22389 7987 22423
rect 9416 22420 9444 22528
rect 9784 22497 9812 22596
rect 10413 22593 10425 22596
rect 10459 22593 10471 22627
rect 10413 22587 10471 22593
rect 10505 22627 10563 22633
rect 10505 22593 10517 22627
rect 10551 22593 10563 22627
rect 10686 22624 10692 22636
rect 10647 22596 10692 22624
rect 10505 22587 10563 22593
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 12406 22624 12434 22664
rect 15473 22661 15485 22695
rect 15519 22692 15531 22695
rect 15654 22692 15660 22704
rect 15519 22664 15660 22692
rect 15519 22661 15531 22664
rect 15473 22655 15531 22661
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 19242 22692 19248 22704
rect 17512 22664 19248 22692
rect 13725 22627 13783 22633
rect 13725 22624 13737 22627
rect 12406 22596 13737 22624
rect 13725 22593 13737 22596
rect 13771 22593 13783 22627
rect 17402 22624 17408 22636
rect 17363 22596 17408 22624
rect 13725 22587 13783 22593
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 17512 22633 17540 22664
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 19613 22695 19671 22701
rect 19613 22661 19625 22695
rect 19659 22692 19671 22695
rect 20346 22692 20352 22704
rect 19659 22664 20352 22692
rect 19659 22661 19671 22664
rect 19613 22655 19671 22661
rect 20346 22652 20352 22664
rect 20404 22652 20410 22704
rect 20441 22695 20499 22701
rect 20441 22661 20453 22695
rect 20487 22692 20499 22695
rect 21266 22692 21272 22704
rect 20487 22664 21272 22692
rect 20487 22661 20499 22664
rect 20441 22655 20499 22661
rect 21266 22652 21272 22664
rect 21324 22692 21330 22704
rect 21361 22695 21419 22701
rect 21361 22692 21373 22695
rect 21324 22664 21373 22692
rect 21324 22652 21330 22664
rect 21361 22661 21373 22664
rect 21407 22692 21419 22695
rect 21818 22692 21824 22704
rect 21407 22664 21824 22692
rect 21407 22661 21419 22664
rect 21361 22655 21419 22661
rect 21818 22652 21824 22664
rect 21876 22652 21882 22704
rect 17497 22627 17555 22633
rect 17497 22593 17509 22627
rect 17543 22593 17555 22627
rect 17497 22587 17555 22593
rect 17586 22584 17592 22636
rect 17644 22624 17650 22636
rect 17773 22627 17831 22633
rect 17644 22596 17689 22624
rect 17644 22584 17650 22596
rect 17773 22593 17785 22627
rect 17819 22593 17831 22627
rect 17773 22587 17831 22593
rect 12250 22556 12256 22568
rect 12211 22528 12256 22556
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 12345 22559 12403 22565
rect 12345 22525 12357 22559
rect 12391 22556 12403 22559
rect 12710 22556 12716 22568
rect 12391 22528 12716 22556
rect 12391 22525 12403 22528
rect 12345 22519 12403 22525
rect 12710 22516 12716 22528
rect 12768 22516 12774 22568
rect 15197 22559 15255 22565
rect 15197 22525 15209 22559
rect 15243 22556 15255 22559
rect 15286 22556 15292 22568
rect 15243 22528 15292 22556
rect 15243 22525 15255 22528
rect 15197 22519 15255 22525
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 15682 22559 15740 22565
rect 15682 22525 15694 22559
rect 15728 22556 15740 22559
rect 15838 22556 15844 22568
rect 15728 22528 15844 22556
rect 15728 22525 15740 22528
rect 15682 22519 15740 22525
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 17788 22556 17816 22587
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 18598 22624 18604 22636
rect 18288 22596 18604 22624
rect 18288 22584 18294 22596
rect 18598 22584 18604 22596
rect 18656 22624 18662 22636
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 18656 22596 18705 22624
rect 18656 22584 18662 22596
rect 18693 22593 18705 22596
rect 18739 22593 18751 22627
rect 19426 22624 19432 22636
rect 19387 22596 19432 22624
rect 18693 22587 18751 22593
rect 19426 22584 19432 22596
rect 19484 22584 19490 22636
rect 20254 22624 20260 22636
rect 20215 22596 20260 22624
rect 20254 22584 20260 22596
rect 20312 22584 20318 22636
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22624 20591 22627
rect 21453 22627 21511 22633
rect 20579 22596 21220 22624
rect 20579 22593 20591 22596
rect 20533 22587 20591 22593
rect 19978 22556 19984 22568
rect 17788 22528 19984 22556
rect 19978 22516 19984 22528
rect 20036 22556 20042 22568
rect 20438 22556 20444 22568
rect 20036 22528 20444 22556
rect 20036 22516 20042 22528
rect 20438 22516 20444 22528
rect 20496 22516 20502 22568
rect 20990 22556 20996 22568
rect 20951 22528 20996 22556
rect 20990 22516 20996 22528
rect 21048 22516 21054 22568
rect 21192 22556 21220 22596
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 21468 22556 21496 22587
rect 21634 22584 21640 22636
rect 21692 22624 21698 22636
rect 22445 22627 22503 22633
rect 22445 22624 22457 22627
rect 21692 22596 22457 22624
rect 21692 22584 21698 22596
rect 22445 22593 22457 22596
rect 22491 22593 22503 22627
rect 22445 22587 22503 22593
rect 21726 22556 21732 22568
rect 21192 22528 21732 22556
rect 21726 22516 21732 22528
rect 21784 22516 21790 22568
rect 22186 22556 22192 22568
rect 22147 22528 22192 22556
rect 22186 22516 22192 22528
rect 22244 22516 22250 22568
rect 9769 22491 9827 22497
rect 9769 22457 9781 22491
rect 9815 22457 9827 22491
rect 9769 22451 9827 22457
rect 10594 22448 10600 22500
rect 10652 22488 10658 22500
rect 11146 22488 11152 22500
rect 10652 22460 10697 22488
rect 10796 22460 11152 22488
rect 10652 22448 10658 22460
rect 10796 22420 10824 22460
rect 11146 22448 11152 22460
rect 11204 22448 11210 22500
rect 11790 22488 11796 22500
rect 11751 22460 11796 22488
rect 11790 22448 11796 22460
rect 11848 22448 11854 22500
rect 12802 22448 12808 22500
rect 12860 22488 12866 22500
rect 13541 22491 13599 22497
rect 13541 22488 13553 22491
rect 12860 22460 13553 22488
rect 12860 22448 12866 22460
rect 13541 22457 13553 22460
rect 13587 22488 13599 22491
rect 14274 22488 14280 22500
rect 13587 22460 14280 22488
rect 13587 22457 13599 22460
rect 13541 22451 13599 22457
rect 14274 22448 14280 22460
rect 14332 22488 14338 22500
rect 18690 22488 18696 22500
rect 14332 22460 18696 22488
rect 14332 22448 14338 22460
rect 18690 22448 18696 22460
rect 18748 22448 18754 22500
rect 9416 22392 10824 22420
rect 7929 22383 7987 22389
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 12529 22423 12587 22429
rect 12529 22420 12541 22423
rect 11112 22392 12541 22420
rect 11112 22380 11118 22392
rect 12529 22389 12541 22392
rect 12575 22389 12587 22423
rect 12529 22383 12587 22389
rect 15746 22380 15752 22432
rect 15804 22420 15810 22432
rect 15841 22423 15899 22429
rect 15841 22420 15853 22423
rect 15804 22392 15853 22420
rect 15804 22380 15810 22392
rect 15841 22389 15853 22392
rect 15887 22389 15899 22423
rect 15841 22383 15899 22389
rect 21177 22423 21235 22429
rect 21177 22389 21189 22423
rect 21223 22420 21235 22423
rect 21542 22420 21548 22432
rect 21223 22392 21548 22420
rect 21223 22389 21235 22392
rect 21177 22383 21235 22389
rect 21542 22380 21548 22392
rect 21600 22380 21606 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 2314 22176 2320 22228
rect 2372 22216 2378 22228
rect 9582 22216 9588 22228
rect 2372 22188 4476 22216
rect 9543 22188 9588 22216
rect 2372 22176 2378 22188
rect 3510 22148 3516 22160
rect 3068 22120 3516 22148
rect 2130 22012 2136 22024
rect 2091 21984 2136 22012
rect 2130 21972 2136 21984
rect 2188 21972 2194 22024
rect 2317 22015 2375 22021
rect 2317 21981 2329 22015
rect 2363 22012 2375 22015
rect 2682 22012 2688 22024
rect 2363 21984 2688 22012
rect 2363 21981 2375 21984
rect 2317 21975 2375 21981
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 2958 22012 2964 22024
rect 2919 21984 2964 22012
rect 2958 21972 2964 21984
rect 3016 21972 3022 22024
rect 3068 22021 3096 22120
rect 3510 22108 3516 22120
rect 3568 22108 3574 22160
rect 4448 22148 4476 22188
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 11701 22219 11759 22225
rect 11701 22185 11713 22219
rect 11747 22216 11759 22219
rect 12250 22216 12256 22228
rect 11747 22188 12256 22216
rect 11747 22185 11759 22188
rect 11701 22179 11759 22185
rect 12250 22176 12256 22188
rect 12308 22176 12314 22228
rect 12710 22216 12716 22228
rect 12671 22188 12716 22216
rect 12710 22176 12716 22188
rect 12768 22176 12774 22228
rect 21361 22219 21419 22225
rect 21361 22185 21373 22219
rect 21407 22216 21419 22219
rect 21634 22216 21640 22228
rect 21407 22188 21640 22216
rect 21407 22185 21419 22188
rect 21361 22179 21419 22185
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 4890 22148 4896 22160
rect 4448 22120 4896 22148
rect 4062 22080 4068 22092
rect 3344 22052 4068 22080
rect 3344 22021 3372 22052
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 21981 3111 22015
rect 3053 21975 3111 21981
rect 3329 22015 3387 22021
rect 3329 21981 3341 22015
rect 3375 21981 3387 22015
rect 3329 21975 3387 21981
rect 3418 21972 3424 22024
rect 3476 22012 3482 22024
rect 4246 22012 4252 22024
rect 3476 21984 3521 22012
rect 4207 21984 4252 22012
rect 3476 21972 3482 21984
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 4448 22021 4476 22120
rect 4890 22108 4896 22120
rect 4948 22108 4954 22160
rect 6086 22108 6092 22160
rect 6144 22148 6150 22160
rect 7834 22148 7840 22160
rect 6144 22120 7840 22148
rect 6144 22108 6150 22120
rect 7834 22108 7840 22120
rect 7892 22108 7898 22160
rect 8294 22148 8300 22160
rect 8255 22120 8300 22148
rect 8294 22108 8300 22120
rect 8352 22108 8358 22160
rect 13265 22151 13323 22157
rect 13265 22117 13277 22151
rect 13311 22148 13323 22151
rect 13311 22120 14320 22148
rect 13311 22117 13323 22120
rect 13265 22111 13323 22117
rect 8938 22080 8944 22092
rect 8496 22052 8944 22080
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 21981 4491 22015
rect 4890 22012 4896 22024
rect 4851 21984 4896 22012
rect 4433 21975 4491 21981
rect 4890 21972 4896 21984
rect 4948 22012 4954 22024
rect 5442 22012 5448 22024
rect 4948 21984 5448 22012
rect 4948 21972 4954 21984
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 8496 22021 8524 22052
rect 8938 22040 8944 22052
rect 8996 22080 9002 22092
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 8996 22052 9873 22080
rect 8996 22040 9002 22052
rect 9861 22049 9873 22052
rect 9907 22049 9919 22083
rect 9861 22043 9919 22049
rect 10045 22083 10103 22089
rect 10045 22049 10057 22083
rect 10091 22080 10103 22083
rect 11054 22080 11060 22092
rect 10091 22052 11060 22080
rect 10091 22049 10103 22052
rect 10045 22043 10103 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 12342 22080 12348 22092
rect 12303 22052 12348 22080
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 14292 22080 14320 22120
rect 17494 22108 17500 22160
rect 17552 22148 17558 22160
rect 17552 22120 19472 22148
rect 17552 22108 17558 22120
rect 16853 22083 16911 22089
rect 14292 22052 14412 22080
rect 8481 22015 8539 22021
rect 8481 21981 8493 22015
rect 8527 21981 8539 22015
rect 8481 21975 8539 21981
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 9582 22012 9588 22024
rect 8619 21984 9588 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 9582 21972 9588 21984
rect 9640 22012 9646 22024
rect 9769 22015 9827 22021
rect 9769 22012 9781 22015
rect 9640 21984 9781 22012
rect 9640 21972 9646 21984
rect 9769 21981 9781 21984
rect 9815 21981 9827 22015
rect 9769 21975 9827 21981
rect 9953 22015 10011 22021
rect 9953 21981 9965 22015
rect 9999 22012 10011 22015
rect 10686 22012 10692 22024
rect 9999 21984 10692 22012
rect 9999 21981 10011 21984
rect 9953 21975 10011 21981
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 11238 21972 11244 22024
rect 11296 22012 11302 22024
rect 11517 22015 11575 22021
rect 11517 22012 11529 22015
rect 11296 21984 11529 22012
rect 11296 21972 11302 21984
rect 11517 21981 11529 21984
rect 11563 21981 11575 22015
rect 11517 21975 11575 21981
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12492 21984 12537 22012
rect 12492 21972 12498 21984
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 12676 21984 13461 22012
rect 12676 21972 12682 21984
rect 13449 21981 13461 21984
rect 13495 21981 13507 22015
rect 13630 22012 13636 22024
rect 13591 21984 13636 22012
rect 13449 21975 13507 21981
rect 13630 21972 13636 21984
rect 13688 21972 13694 22024
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 21981 13783 22015
rect 14274 22012 14280 22024
rect 14235 21984 14280 22012
rect 13725 21975 13783 21981
rect 2225 21947 2283 21953
rect 2225 21913 2237 21947
rect 2271 21944 2283 21947
rect 2976 21944 3004 21972
rect 2271 21916 3004 21944
rect 3145 21947 3203 21953
rect 2271 21913 2283 21916
rect 2225 21907 2283 21913
rect 3145 21913 3157 21947
rect 3191 21944 3203 21947
rect 3602 21944 3608 21956
rect 3191 21916 3608 21944
rect 3191 21913 3203 21916
rect 3145 21907 3203 21913
rect 3602 21904 3608 21916
rect 3660 21904 3666 21956
rect 4341 21947 4399 21953
rect 4341 21913 4353 21947
rect 4387 21944 4399 21947
rect 5138 21947 5196 21953
rect 5138 21944 5150 21947
rect 4387 21916 5150 21944
rect 4387 21913 4399 21916
rect 4341 21907 4399 21913
rect 5138 21913 5150 21916
rect 5184 21913 5196 21947
rect 5138 21907 5196 21913
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 8297 21947 8355 21953
rect 5684 21916 6776 21944
rect 5684 21904 5690 21916
rect 2777 21879 2835 21885
rect 2777 21845 2789 21879
rect 2823 21876 2835 21879
rect 3234 21876 3240 21888
rect 2823 21848 3240 21876
rect 2823 21845 2835 21848
rect 2777 21839 2835 21845
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 6273 21879 6331 21885
rect 6273 21845 6285 21879
rect 6319 21876 6331 21879
rect 6638 21876 6644 21888
rect 6319 21848 6644 21876
rect 6319 21845 6331 21848
rect 6273 21839 6331 21845
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 6748 21876 6776 21916
rect 8297 21913 8309 21947
rect 8343 21944 8355 21947
rect 9398 21944 9404 21956
rect 8343 21916 9404 21944
rect 8343 21913 8355 21916
rect 8297 21907 8355 21913
rect 9398 21904 9404 21916
rect 9456 21904 9462 21956
rect 11054 21904 11060 21956
rect 11112 21944 11118 21956
rect 11149 21947 11207 21953
rect 11149 21944 11161 21947
rect 11112 21916 11161 21944
rect 11112 21904 11118 21916
rect 11149 21913 11161 21916
rect 11195 21913 11207 21947
rect 11149 21907 11207 21913
rect 11425 21947 11483 21953
rect 11425 21913 11437 21947
rect 11471 21944 11483 21947
rect 11882 21944 11888 21956
rect 11471 21916 11888 21944
rect 11471 21913 11483 21916
rect 11425 21907 11483 21913
rect 11882 21904 11888 21916
rect 11940 21904 11946 21956
rect 13740 21944 13768 21975
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 14384 22012 14412 22052
rect 16853 22049 16865 22083
rect 16899 22080 16911 22083
rect 17218 22080 17224 22092
rect 16899 22052 17224 22080
rect 16899 22049 16911 22052
rect 16853 22043 16911 22049
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 17862 22040 17868 22092
rect 17920 22080 17926 22092
rect 17920 22052 18920 22080
rect 17920 22040 17926 22052
rect 14533 22015 14591 22021
rect 14533 22012 14545 22015
rect 14384 21984 14545 22012
rect 14533 21981 14545 21984
rect 14579 21981 14591 22015
rect 14533 21975 14591 21981
rect 15378 21972 15384 22024
rect 15436 22012 15442 22024
rect 16482 22012 16488 22024
rect 15436 21984 16488 22012
rect 15436 21972 15442 21984
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 16945 22015 17003 22021
rect 16945 21981 16957 22015
rect 16991 22012 17003 22015
rect 17034 22012 17040 22024
rect 16991 21984 17040 22012
rect 16991 21981 17003 21984
rect 16945 21975 17003 21981
rect 17034 21972 17040 21984
rect 17092 21972 17098 22024
rect 17586 21972 17592 22024
rect 17644 22012 17650 22024
rect 17957 22015 18015 22021
rect 17957 22012 17969 22015
rect 17644 21984 17969 22012
rect 17644 21972 17650 21984
rect 17957 21981 17969 21984
rect 18003 21981 18015 22015
rect 17957 21975 18015 21981
rect 18049 22015 18107 22021
rect 18049 21981 18061 22015
rect 18095 22012 18107 22015
rect 18506 22012 18512 22024
rect 18095 21984 18512 22012
rect 18095 21981 18107 21984
rect 18049 21975 18107 21981
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 18690 22012 18696 22024
rect 18651 21984 18696 22012
rect 18690 21972 18696 21984
rect 18748 21972 18754 22024
rect 18892 22021 18920 22052
rect 19444 22021 19472 22120
rect 22649 22083 22707 22089
rect 22649 22080 22661 22083
rect 21744 22052 22661 22080
rect 21744 22024 21772 22052
rect 22649 22049 22661 22052
rect 22695 22049 22707 22083
rect 22649 22043 22707 22049
rect 18877 22015 18935 22021
rect 18877 21981 18889 22015
rect 18923 21981 18935 22015
rect 18877 21975 18935 21981
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 22012 19487 22015
rect 19978 22012 19984 22024
rect 19475 21984 19984 22012
rect 19475 21981 19487 21984
rect 19429 21975 19487 21981
rect 19978 21972 19984 21984
rect 20036 21972 20042 22024
rect 21542 22012 21548 22024
rect 21503 21984 21548 22012
rect 21542 21972 21548 21984
rect 21600 21972 21606 22024
rect 21726 22012 21732 22024
rect 21687 21984 21732 22012
rect 21726 21972 21732 21984
rect 21784 21972 21790 22024
rect 21818 21972 21824 22024
rect 21876 22012 21882 22024
rect 22373 22015 22431 22021
rect 21876 21984 21921 22012
rect 21876 21972 21882 21984
rect 22373 21981 22385 22015
rect 22419 22012 22431 22015
rect 23198 22012 23204 22024
rect 22419 21984 23204 22012
rect 22419 21981 22431 21984
rect 22373 21975 22431 21981
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 13906 21944 13912 21956
rect 13740 21916 13912 21944
rect 13906 21904 13912 21916
rect 13964 21944 13970 21956
rect 15746 21944 15752 21956
rect 13964 21916 15752 21944
rect 13964 21904 13970 21916
rect 15746 21904 15752 21916
rect 15804 21904 15810 21956
rect 15930 21904 15936 21956
rect 15988 21944 15994 21956
rect 17773 21947 17831 21953
rect 17773 21944 17785 21947
rect 15988 21916 17785 21944
rect 15988 21904 15994 21916
rect 17773 21913 17785 21916
rect 17819 21913 17831 21947
rect 17773 21907 17831 21913
rect 18785 21947 18843 21953
rect 18785 21913 18797 21947
rect 18831 21944 18843 21947
rect 19674 21947 19732 21953
rect 19674 21944 19686 21947
rect 18831 21916 19686 21944
rect 18831 21913 18843 21916
rect 18785 21907 18843 21913
rect 19674 21913 19686 21916
rect 19720 21913 19732 21947
rect 19674 21907 19732 21913
rect 9858 21876 9864 21888
rect 6748 21848 9864 21876
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 11330 21876 11336 21888
rect 11291 21848 11336 21876
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 15194 21836 15200 21888
rect 15252 21876 15258 21888
rect 15657 21879 15715 21885
rect 15657 21876 15669 21879
rect 15252 21848 15669 21876
rect 15252 21836 15258 21848
rect 15657 21845 15669 21848
rect 15703 21845 15715 21879
rect 15657 21839 15715 21845
rect 17034 21836 17040 21888
rect 17092 21876 17098 21888
rect 17313 21879 17371 21885
rect 17313 21876 17325 21879
rect 17092 21848 17325 21876
rect 17092 21836 17098 21848
rect 17313 21845 17325 21848
rect 17359 21845 17371 21879
rect 17313 21839 17371 21845
rect 17402 21836 17408 21888
rect 17460 21876 17466 21888
rect 17871 21879 17929 21885
rect 17871 21876 17883 21879
rect 17460 21848 17883 21876
rect 17460 21836 17466 21848
rect 17871 21845 17883 21848
rect 17917 21845 17929 21879
rect 17871 21839 17929 21845
rect 20162 21836 20168 21888
rect 20220 21876 20226 21888
rect 20809 21879 20867 21885
rect 20809 21876 20821 21879
rect 20220 21848 20821 21876
rect 20220 21836 20226 21848
rect 20809 21845 20821 21848
rect 20855 21845 20867 21879
rect 20809 21839 20867 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2774 21632 2780 21684
rect 2832 21672 2838 21684
rect 2832 21644 2877 21672
rect 2832 21632 2838 21644
rect 4246 21632 4252 21684
rect 4304 21672 4310 21684
rect 4341 21675 4399 21681
rect 4341 21672 4353 21675
rect 4304 21644 4353 21672
rect 4304 21632 4310 21644
rect 4341 21641 4353 21644
rect 4387 21641 4399 21675
rect 7374 21672 7380 21684
rect 7335 21644 7380 21672
rect 4341 21635 4399 21641
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 7484 21644 8984 21672
rect 2130 21564 2136 21616
rect 2188 21604 2194 21616
rect 2409 21607 2467 21613
rect 2409 21604 2421 21607
rect 2188 21576 2421 21604
rect 2188 21564 2194 21576
rect 2409 21573 2421 21576
rect 2455 21604 2467 21607
rect 4982 21604 4988 21616
rect 2455 21576 4988 21604
rect 2455 21573 2467 21576
rect 2409 21567 2467 21573
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21505 2651 21539
rect 2593 21499 2651 21505
rect 2608 21468 2636 21499
rect 2866 21496 2872 21548
rect 2924 21536 2930 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 2924 21508 3433 21536
rect 2924 21496 2930 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 4525 21539 4583 21545
rect 4525 21536 4537 21539
rect 3421 21499 3479 21505
rect 3804 21508 4537 21536
rect 3050 21468 3056 21480
rect 2608 21440 3056 21468
rect 3050 21428 3056 21440
rect 3108 21428 3114 21480
rect 3326 21468 3332 21480
rect 3287 21440 3332 21468
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 3804 21409 3832 21508
rect 4525 21505 4537 21508
rect 4571 21505 4583 21539
rect 4525 21499 4583 21505
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21536 4675 21539
rect 4706 21536 4712 21548
rect 4663 21508 4712 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 4706 21496 4712 21508
rect 4764 21496 4770 21548
rect 4908 21545 4936 21576
rect 4982 21564 4988 21576
rect 5040 21604 5046 21616
rect 6733 21607 6791 21613
rect 6733 21604 6745 21607
rect 5040 21576 6745 21604
rect 5040 21564 5046 21576
rect 6733 21573 6745 21576
rect 6779 21604 6791 21607
rect 7484 21604 7512 21644
rect 8956 21604 8984 21644
rect 9582 21632 9588 21684
rect 9640 21672 9646 21684
rect 9769 21675 9827 21681
rect 9769 21672 9781 21675
rect 9640 21644 9781 21672
rect 9640 21632 9646 21644
rect 9769 21641 9781 21644
rect 9815 21641 9827 21675
rect 9769 21635 9827 21641
rect 9858 21632 9864 21684
rect 9916 21672 9922 21684
rect 12526 21672 12532 21684
rect 9916 21644 12532 21672
rect 9916 21632 9922 21644
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 13630 21632 13636 21684
rect 13688 21672 13694 21684
rect 14921 21675 14979 21681
rect 14921 21672 14933 21675
rect 13688 21644 14933 21672
rect 13688 21632 13694 21644
rect 14921 21641 14933 21644
rect 14967 21641 14979 21675
rect 14921 21635 14979 21641
rect 15396 21644 15608 21672
rect 11974 21604 11980 21616
rect 6779 21576 7512 21604
rect 7576 21576 8892 21604
rect 8956 21576 11980 21604
rect 6779 21573 6791 21576
rect 6733 21567 6791 21573
rect 4893 21539 4951 21545
rect 4893 21505 4905 21539
rect 4939 21505 4951 21539
rect 5626 21536 5632 21548
rect 5587 21508 5632 21536
rect 4893 21499 4951 21505
rect 5626 21496 5632 21508
rect 5684 21496 5690 21548
rect 6638 21536 6644 21548
rect 6599 21508 6644 21536
rect 6638 21496 6644 21508
rect 6696 21496 6702 21548
rect 7576 21545 7604 21576
rect 8864 21548 8892 21576
rect 11974 21564 11980 21576
rect 12032 21564 12038 21616
rect 15396 21604 15424 21644
rect 12406 21576 15424 21604
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21505 7619 21539
rect 7834 21536 7840 21548
rect 7795 21508 7840 21536
rect 7561 21499 7619 21505
rect 7834 21496 7840 21508
rect 7892 21496 7898 21548
rect 8386 21536 8392 21548
rect 8347 21508 8392 21536
rect 8386 21496 8392 21508
rect 8444 21496 8450 21548
rect 8570 21536 8576 21548
rect 8531 21508 8576 21536
rect 8570 21496 8576 21508
rect 8628 21496 8634 21548
rect 8662 21496 8668 21548
rect 8720 21536 8726 21548
rect 8846 21536 8852 21548
rect 8720 21508 8765 21536
rect 8807 21508 8852 21536
rect 8720 21496 8726 21508
rect 8846 21496 8852 21508
rect 8904 21496 8910 21548
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 9585 21539 9643 21545
rect 8996 21508 9041 21536
rect 8996 21496 9002 21508
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9858 21536 9864 21548
rect 9631 21508 9864 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9858 21496 9864 21508
rect 9916 21496 9922 21548
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21536 10747 21539
rect 10870 21536 10876 21548
rect 10735 21508 10876 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21536 11023 21539
rect 11790 21536 11796 21548
rect 11011 21508 11796 21536
rect 11011 21505 11023 21508
rect 10965 21499 11023 21505
rect 11790 21496 11796 21508
rect 11848 21496 11854 21548
rect 12253 21539 12311 21545
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 12406 21536 12434 21576
rect 15470 21564 15476 21616
rect 15528 21564 15534 21616
rect 15580 21604 15608 21644
rect 15654 21632 15660 21684
rect 15712 21672 15718 21684
rect 17402 21672 17408 21684
rect 15712 21644 17408 21672
rect 15712 21632 15718 21644
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 17862 21632 17868 21684
rect 17920 21672 17926 21684
rect 19797 21675 19855 21681
rect 19797 21672 19809 21675
rect 17920 21644 19809 21672
rect 17920 21632 17926 21644
rect 19797 21641 19809 21644
rect 19843 21641 19855 21675
rect 19797 21635 19855 21641
rect 21085 21675 21143 21681
rect 21085 21641 21097 21675
rect 21131 21672 21143 21675
rect 22002 21672 22008 21684
rect 21131 21644 22008 21672
rect 21131 21641 21143 21644
rect 21085 21635 21143 21641
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 23198 21632 23204 21684
rect 23256 21672 23262 21684
rect 23845 21675 23903 21681
rect 23845 21672 23857 21675
rect 23256 21644 23857 21672
rect 23256 21632 23262 21644
rect 23845 21641 23857 21644
rect 23891 21641 23903 21675
rect 23845 21635 23903 21641
rect 19426 21604 19432 21616
rect 15580 21576 19432 21604
rect 19426 21564 19432 21576
rect 19484 21604 19490 21616
rect 20162 21604 20168 21616
rect 19484 21576 20168 21604
rect 19484 21564 19490 21576
rect 15194 21536 15200 21548
rect 12299 21508 12434 21536
rect 15155 21508 15200 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 15488 21536 15516 21564
rect 15657 21539 15715 21545
rect 15657 21536 15669 21539
rect 15488 21508 15669 21536
rect 15657 21505 15669 21508
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 16942 21496 16948 21548
rect 17000 21536 17006 21548
rect 17129 21539 17187 21545
rect 17129 21536 17141 21539
rect 17000 21508 17141 21536
rect 17000 21496 17006 21508
rect 17129 21505 17141 21508
rect 17175 21505 17187 21539
rect 17129 21499 17187 21505
rect 17396 21539 17454 21545
rect 17396 21505 17408 21539
rect 17442 21536 17454 21539
rect 17678 21536 17684 21548
rect 17442 21508 17684 21536
rect 17442 21505 17454 21508
rect 17396 21499 17454 21505
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 19536 21545 19564 21576
rect 20162 21564 20168 21576
rect 20220 21564 20226 21616
rect 20809 21607 20867 21613
rect 20809 21573 20821 21607
rect 20855 21604 20867 21607
rect 20898 21604 20904 21616
rect 20855 21576 20904 21604
rect 20855 21573 20867 21576
rect 20809 21567 20867 21573
rect 20898 21564 20904 21576
rect 20956 21564 20962 21616
rect 20993 21607 21051 21613
rect 20993 21573 21005 21607
rect 21039 21604 21051 21607
rect 21726 21604 21732 21616
rect 21039 21576 21732 21604
rect 21039 21573 21051 21576
rect 20993 21567 21051 21573
rect 21726 21564 21732 21576
rect 21784 21564 21790 21616
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 19610 21496 19616 21548
rect 19668 21536 19674 21548
rect 20530 21536 20536 21548
rect 19668 21508 20536 21536
rect 19668 21496 19674 21508
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 21818 21536 21824 21548
rect 21131 21508 21824 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22732 21539 22790 21545
rect 22732 21505 22744 21539
rect 22778 21536 22790 21539
rect 23014 21536 23020 21548
rect 22778 21508 23020 21536
rect 22778 21505 22790 21508
rect 22732 21499 22790 21505
rect 23014 21496 23020 21508
rect 23072 21496 23078 21548
rect 4798 21468 4804 21480
rect 4759 21440 4804 21468
rect 4798 21428 4804 21440
rect 4856 21428 4862 21480
rect 5721 21471 5779 21477
rect 5721 21437 5733 21471
rect 5767 21468 5779 21471
rect 6086 21468 6092 21480
rect 5767 21440 6092 21468
rect 5767 21437 5779 21440
rect 5721 21431 5779 21437
rect 6086 21428 6092 21440
rect 6144 21428 6150 21480
rect 3789 21403 3847 21409
rect 3789 21369 3801 21403
rect 3835 21369 3847 21403
rect 5994 21400 6000 21412
rect 5955 21372 6000 21400
rect 3789 21363 3847 21369
rect 5994 21360 6000 21372
rect 6052 21360 6058 21412
rect 6656 21332 6684 21496
rect 7374 21428 7380 21480
rect 7432 21468 7438 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7432 21440 7665 21468
rect 7432 21428 7438 21440
rect 7653 21437 7665 21440
rect 7699 21468 7711 21471
rect 8956 21468 8984 21496
rect 7699 21440 8984 21468
rect 7699 21437 7711 21440
rect 7653 21431 7711 21437
rect 9306 21428 9312 21480
rect 9364 21468 9370 21480
rect 9401 21471 9459 21477
rect 9401 21468 9413 21471
rect 9364 21440 9413 21468
rect 9364 21428 9370 21440
rect 9401 21437 9413 21440
rect 9447 21437 9459 21471
rect 10778 21468 10784 21480
rect 10739 21440 10784 21468
rect 9401 21431 9459 21437
rect 10778 21428 10784 21440
rect 10836 21428 10842 21480
rect 12161 21471 12219 21477
rect 12161 21468 12173 21471
rect 10888 21440 12173 21468
rect 7745 21403 7803 21409
rect 7745 21369 7757 21403
rect 7791 21400 7803 21403
rect 7926 21400 7932 21412
rect 7791 21372 7932 21400
rect 7791 21369 7803 21372
rect 7745 21363 7803 21369
rect 7926 21360 7932 21372
rect 7984 21360 7990 21412
rect 8128 21372 8524 21400
rect 8128 21332 8156 21372
rect 8496 21344 8524 21372
rect 8846 21360 8852 21412
rect 8904 21400 8910 21412
rect 9324 21400 9352 21428
rect 8904 21372 9352 21400
rect 8904 21360 8910 21372
rect 6656 21304 8156 21332
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 10888 21332 10916 21440
rect 12161 21437 12173 21440
rect 12207 21468 12219 21471
rect 12526 21468 12532 21480
rect 12207 21440 12532 21468
rect 12207 21437 12219 21440
rect 12161 21431 12219 21437
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 15473 21471 15531 21477
rect 15473 21437 15485 21471
rect 15519 21468 15531 21471
rect 17034 21468 17040 21480
rect 15519 21440 17040 21468
rect 15519 21437 15531 21440
rect 15473 21431 15531 21437
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 19978 21428 19984 21480
rect 20036 21468 20042 21480
rect 22186 21468 22192 21480
rect 20036 21440 22192 21468
rect 20036 21428 20042 21440
rect 22186 21428 22192 21440
rect 22244 21468 22250 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22244 21440 22477 21468
rect 22244 21428 22250 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 11330 21400 11336 21412
rect 10980 21372 11336 21400
rect 10980 21341 11008 21372
rect 11330 21360 11336 21372
rect 11388 21400 11394 21412
rect 12621 21403 12679 21409
rect 12621 21400 12633 21403
rect 11388 21372 12633 21400
rect 11388 21360 11394 21372
rect 12621 21369 12633 21372
rect 12667 21369 12679 21403
rect 12621 21363 12679 21369
rect 8536 21304 10916 21332
rect 10965 21335 11023 21341
rect 8536 21292 8542 21304
rect 10965 21301 10977 21335
rect 11011 21301 11023 21335
rect 11146 21332 11152 21344
rect 11107 21304 11152 21332
rect 10965 21295 11023 21301
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 15286 21332 15292 21344
rect 15247 21304 15292 21332
rect 15286 21292 15292 21304
rect 15344 21292 15350 21344
rect 15378 21292 15384 21344
rect 15436 21332 15442 21344
rect 15436 21304 15481 21332
rect 15436 21292 15442 21304
rect 16758 21292 16764 21344
rect 16816 21332 16822 21344
rect 18509 21335 18567 21341
rect 18509 21332 18521 21335
rect 16816 21304 18521 21332
rect 16816 21292 16822 21304
rect 18509 21301 18521 21304
rect 18555 21301 18567 21335
rect 18509 21295 18567 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 6730 21128 6736 21140
rect 2516 21100 6736 21128
rect 2317 21063 2375 21069
rect 2317 21029 2329 21063
rect 2363 21029 2375 21063
rect 2317 21023 2375 21029
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 2332 20924 2360 21023
rect 2516 20933 2544 21100
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 6825 21131 6883 21137
rect 6825 21097 6837 21131
rect 6871 21097 6883 21131
rect 7098 21128 7104 21140
rect 7059 21100 7104 21128
rect 6825 21091 6883 21097
rect 5813 21063 5871 21069
rect 5813 21029 5825 21063
rect 5859 21060 5871 21063
rect 6270 21060 6276 21072
rect 5859 21032 6276 21060
rect 5859 21029 5871 21032
rect 5813 21023 5871 21029
rect 6270 21020 6276 21032
rect 6328 21020 6334 21072
rect 6840 21060 6868 21091
rect 7098 21088 7104 21100
rect 7156 21088 7162 21140
rect 7926 21128 7932 21140
rect 7887 21100 7932 21128
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 8570 21128 8576 21140
rect 8220 21100 8576 21128
rect 7006 21060 7012 21072
rect 6840 21032 7012 21060
rect 7006 21020 7012 21032
rect 7064 21020 7070 21072
rect 8220 21060 8248 21100
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 9398 21088 9404 21140
rect 9456 21128 9462 21140
rect 9585 21131 9643 21137
rect 9585 21128 9597 21131
rect 9456 21100 9597 21128
rect 9456 21088 9462 21100
rect 9585 21097 9597 21100
rect 9631 21097 9643 21131
rect 9585 21091 9643 21097
rect 10413 21131 10471 21137
rect 10413 21097 10425 21131
rect 10459 21128 10471 21131
rect 10594 21128 10600 21140
rect 10459 21100 10600 21128
rect 10459 21097 10471 21100
rect 10413 21091 10471 21097
rect 10594 21088 10600 21100
rect 10652 21088 10658 21140
rect 10781 21131 10839 21137
rect 10781 21097 10793 21131
rect 10827 21128 10839 21131
rect 11146 21128 11152 21140
rect 10827 21100 11152 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 12250 21128 12256 21140
rect 11256 21100 12256 21128
rect 7760 21032 8248 21060
rect 4246 20992 4252 21004
rect 3252 20964 4252 20992
rect 3252 20936 3280 20964
rect 4246 20952 4252 20964
rect 4304 20952 4310 21004
rect 5537 20995 5595 21001
rect 5537 20961 5549 20995
rect 5583 20992 5595 20995
rect 6825 20995 6883 21001
rect 6825 20992 6837 20995
rect 5583 20964 6837 20992
rect 5583 20961 5595 20964
rect 5537 20955 5595 20961
rect 6825 20961 6837 20964
rect 6871 20961 6883 20995
rect 6825 20955 6883 20961
rect 1627 20896 2360 20924
rect 2501 20927 2559 20933
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 2501 20893 2513 20927
rect 2547 20893 2559 20927
rect 3234 20924 3240 20936
rect 3195 20896 3240 20924
rect 2501 20887 2559 20893
rect 3234 20884 3240 20896
rect 3292 20884 3298 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20924 3479 20927
rect 3970 20924 3976 20936
rect 3467 20896 3976 20924
rect 3467 20893 3479 20896
rect 3421 20887 3479 20893
rect 3970 20884 3976 20896
rect 4028 20884 4034 20936
rect 5626 20884 5632 20936
rect 5684 20924 5690 20936
rect 5721 20927 5779 20933
rect 5721 20924 5733 20927
rect 5684 20896 5733 20924
rect 5684 20884 5690 20896
rect 5721 20893 5733 20896
rect 5767 20893 5779 20927
rect 5902 20924 5908 20936
rect 5863 20896 5908 20924
rect 5721 20887 5779 20893
rect 5902 20884 5908 20896
rect 5960 20884 5966 20936
rect 5994 20884 6000 20936
rect 6052 20924 6058 20936
rect 6362 20924 6368 20936
rect 6052 20896 6368 20924
rect 6052 20884 6058 20896
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 6546 20924 6552 20936
rect 6507 20896 6552 20924
rect 6546 20884 6552 20896
rect 6604 20884 6610 20936
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7760 20924 7788 21032
rect 8294 21020 8300 21072
rect 8352 21060 8358 21072
rect 10689 21063 10747 21069
rect 10689 21060 10701 21063
rect 8352 21032 10701 21060
rect 8352 21020 8358 21032
rect 10689 21029 10701 21032
rect 10735 21029 10747 21063
rect 11256 21060 11284 21100
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 13449 21131 13507 21137
rect 13449 21128 13461 21131
rect 12492 21100 13461 21128
rect 12492 21088 12498 21100
rect 13449 21097 13461 21100
rect 13495 21097 13507 21131
rect 13449 21091 13507 21097
rect 12345 21063 12403 21069
rect 12345 21060 12357 21063
rect 10689 21023 10747 21029
rect 10796 21032 11284 21060
rect 11716 21032 12357 21060
rect 7834 20952 7840 21004
rect 7892 20992 7898 21004
rect 9217 20995 9275 21001
rect 9217 20992 9229 20995
rect 7892 20964 9229 20992
rect 7892 20952 7898 20964
rect 9217 20961 9229 20964
rect 9263 20961 9275 20995
rect 9217 20955 9275 20961
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 10796 20992 10824 21032
rect 9732 20964 10824 20992
rect 10873 20995 10931 21001
rect 9732 20952 9738 20964
rect 10873 20961 10885 20995
rect 10919 20992 10931 20995
rect 11514 20992 11520 21004
rect 10919 20964 11520 20992
rect 10919 20961 10931 20964
rect 10873 20955 10931 20961
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 11716 20936 11744 21032
rect 12345 21029 12357 21032
rect 12391 21029 12403 21063
rect 13464 21060 13492 21091
rect 15286 21088 15292 21140
rect 15344 21128 15350 21140
rect 15381 21131 15439 21137
rect 15381 21128 15393 21131
rect 15344 21100 15393 21128
rect 15344 21088 15350 21100
rect 15381 21097 15393 21100
rect 15427 21097 15439 21131
rect 15381 21091 15439 21097
rect 15838 21088 15844 21140
rect 15896 21128 15902 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 15896 21100 16681 21128
rect 15896 21088 15902 21100
rect 16669 21097 16681 21100
rect 16715 21097 16727 21131
rect 17678 21128 17684 21140
rect 17639 21100 17684 21128
rect 16669 21091 16727 21097
rect 17678 21088 17684 21100
rect 17736 21088 17742 21140
rect 18690 21088 18696 21140
rect 18748 21128 18754 21140
rect 19705 21131 19763 21137
rect 19705 21128 19717 21131
rect 18748 21100 19717 21128
rect 18748 21088 18754 21100
rect 19705 21097 19717 21100
rect 19751 21097 19763 21131
rect 19705 21091 19763 21097
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 21266 21128 21272 21140
rect 21048 21100 21272 21128
rect 21048 21088 21054 21100
rect 21266 21088 21272 21100
rect 21324 21128 21330 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 21324 21100 21465 21128
rect 21324 21088 21330 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 23014 21128 23020 21140
rect 22975 21100 23020 21128
rect 21453 21091 21511 21097
rect 23014 21088 23020 21100
rect 23072 21088 23078 21140
rect 17494 21060 17500 21072
rect 13464 21032 17500 21060
rect 12345 21023 12403 21029
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 18506 21060 18512 21072
rect 17788 21032 18512 21060
rect 11882 20992 11888 21004
rect 11843 20964 11888 20992
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 14642 20992 14648 21004
rect 13372 20964 14648 20992
rect 8113 20927 8171 20933
rect 8113 20924 8125 20927
rect 6972 20896 8125 20924
rect 6972 20884 6978 20896
rect 8113 20893 8125 20896
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 8297 20927 8355 20933
rect 8297 20893 8309 20927
rect 8343 20893 8355 20927
rect 8297 20887 8355 20893
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 8478 20924 8484 20936
rect 8435 20896 8484 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 2958 20816 2964 20868
rect 3016 20856 3022 20868
rect 4433 20859 4491 20865
rect 4433 20856 4445 20859
rect 3016 20828 4445 20856
rect 3016 20816 3022 20828
rect 4433 20825 4445 20828
rect 4479 20825 4491 20859
rect 4433 20819 4491 20825
rect 4617 20859 4675 20865
rect 4617 20825 4629 20859
rect 4663 20856 4675 20859
rect 6086 20856 6092 20868
rect 4663 20828 6092 20856
rect 4663 20825 4675 20828
rect 4617 20819 4675 20825
rect 6086 20816 6092 20828
rect 6144 20856 6150 20868
rect 8312 20856 8340 20887
rect 8478 20884 8484 20896
rect 8536 20884 8542 20936
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20924 9367 20927
rect 10594 20924 10600 20936
rect 9355 20896 10600 20924
rect 9355 20893 9367 20896
rect 9309 20887 9367 20893
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 10962 20924 10968 20936
rect 10923 20896 10968 20924
rect 10962 20884 10968 20896
rect 11020 20884 11026 20936
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20924 11207 20927
rect 11238 20924 11244 20936
rect 11195 20896 11244 20924
rect 11195 20893 11207 20896
rect 11149 20887 11207 20893
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20893 11667 20927
rect 11609 20887 11667 20893
rect 8662 20856 8668 20868
rect 6144 20828 8668 20856
rect 6144 20816 6150 20828
rect 8662 20816 8668 20828
rect 8720 20856 8726 20868
rect 9674 20856 9680 20868
rect 8720 20828 9680 20856
rect 8720 20816 8726 20828
rect 9674 20816 9680 20828
rect 9732 20816 9738 20868
rect 11054 20816 11060 20868
rect 11112 20856 11118 20868
rect 11624 20856 11652 20887
rect 11698 20884 11704 20936
rect 11756 20924 11762 20936
rect 12342 20924 12348 20936
rect 11756 20896 11801 20924
rect 12303 20896 12348 20924
rect 11756 20884 11762 20896
rect 12342 20884 12348 20896
rect 12400 20884 12406 20936
rect 12526 20924 12532 20936
rect 12487 20896 12532 20924
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 13372 20865 13400 20964
rect 14642 20952 14648 20964
rect 14700 20992 14706 21004
rect 16758 20992 16764 21004
rect 14700 20964 16764 20992
rect 14700 20952 14706 20964
rect 16758 20952 16764 20964
rect 16816 20952 16822 21004
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 15654 20924 15660 20936
rect 15611 20896 15660 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 15838 20924 15844 20936
rect 15799 20896 15844 20924
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 17788 20924 17816 21032
rect 18506 21020 18512 21032
rect 18564 21020 18570 21072
rect 19610 21060 19616 21072
rect 19571 21032 19616 21060
rect 19610 21020 19616 21032
rect 19668 21020 19674 21072
rect 20254 21060 20260 21072
rect 19720 21032 20260 21060
rect 18601 20995 18659 21001
rect 18601 20992 18613 20995
rect 17972 20964 18613 20992
rect 16316 20896 17816 20924
rect 13357 20859 13415 20865
rect 13357 20856 13369 20859
rect 11112 20828 13369 20856
rect 11112 20816 11118 20828
rect 13357 20825 13369 20828
rect 13403 20825 13415 20859
rect 13357 20819 13415 20825
rect 15749 20859 15807 20865
rect 15749 20825 15761 20859
rect 15795 20856 15807 20859
rect 15930 20856 15936 20868
rect 15795 20828 15936 20856
rect 15795 20825 15807 20828
rect 15749 20819 15807 20825
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 16316 20865 16344 20896
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 17972 20933 18000 20964
rect 18601 20961 18613 20964
rect 18647 20961 18659 20995
rect 18601 20955 18659 20961
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20992 18843 20995
rect 18966 20992 18972 21004
rect 18831 20964 18972 20992
rect 18831 20961 18843 20964
rect 18785 20955 18843 20961
rect 18966 20952 18972 20964
rect 19024 20992 19030 21004
rect 19720 20992 19748 21032
rect 20254 21020 20260 21032
rect 20312 21020 20318 21072
rect 22186 21020 22192 21072
rect 22244 21060 22250 21072
rect 22373 21063 22431 21069
rect 22373 21060 22385 21063
rect 22244 21032 22385 21060
rect 22244 21020 22250 21032
rect 22373 21029 22385 21032
rect 22419 21029 22431 21063
rect 22373 21023 22431 21029
rect 19024 20964 19748 20992
rect 19797 20995 19855 21001
rect 19024 20952 19030 20964
rect 19797 20961 19809 20995
rect 19843 20992 19855 20995
rect 20438 20992 20444 21004
rect 19843 20964 20444 20992
rect 19843 20961 19855 20964
rect 19797 20955 19855 20961
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 22097 20995 22155 21001
rect 22097 20992 22109 20995
rect 21784 20964 22109 20992
rect 21784 20952 21790 20964
rect 22097 20961 22109 20964
rect 22143 20961 22155 20995
rect 22097 20955 22155 20961
rect 22557 20995 22615 21001
rect 22557 20961 22569 20995
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 17957 20927 18015 20933
rect 17957 20924 17969 20927
rect 17920 20896 17969 20924
rect 17920 20884 17926 20896
rect 17957 20893 17969 20896
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 18322 20884 18328 20936
rect 18380 20924 18386 20936
rect 18509 20927 18567 20933
rect 18509 20924 18521 20927
rect 18380 20896 18521 20924
rect 18380 20884 18386 20896
rect 18509 20893 18521 20896
rect 18555 20924 18567 20927
rect 19242 20924 19248 20936
rect 18555 20896 19248 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 20162 20924 20168 20936
rect 19567 20896 20168 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 20162 20884 20168 20896
rect 20220 20924 20226 20936
rect 20346 20924 20352 20936
rect 20220 20896 20352 20924
rect 20220 20884 20226 20896
rect 20346 20884 20352 20896
rect 20404 20924 20410 20936
rect 20898 20924 20904 20936
rect 20404 20896 20904 20924
rect 20404 20884 20410 20896
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 21082 20924 21088 20936
rect 21043 20896 21088 20924
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 22572 20924 22600 20955
rect 23201 20927 23259 20933
rect 23201 20924 23213 20927
rect 22572 20896 23213 20924
rect 23201 20893 23213 20896
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 16301 20859 16359 20865
rect 16301 20825 16313 20859
rect 16347 20825 16359 20859
rect 16301 20819 16359 20825
rect 16485 20859 16543 20865
rect 16485 20825 16497 20859
rect 16531 20856 16543 20859
rect 17586 20856 17592 20868
rect 16531 20828 17592 20856
rect 16531 20825 16543 20828
rect 16485 20819 16543 20825
rect 1762 20788 1768 20800
rect 1723 20760 1768 20788
rect 1762 20748 1768 20760
rect 1820 20748 1826 20800
rect 3418 20788 3424 20800
rect 3379 20760 3424 20788
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 7006 20748 7012 20800
rect 7064 20788 7070 20800
rect 9766 20788 9772 20800
rect 7064 20760 9772 20788
rect 7064 20748 7070 20760
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 11885 20791 11943 20797
rect 11885 20757 11897 20791
rect 11931 20788 11943 20791
rect 12158 20788 12164 20800
rect 11931 20760 12164 20788
rect 11931 20757 11943 20760
rect 11885 20751 11943 20757
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 15102 20748 15108 20800
rect 15160 20788 15166 20800
rect 16500 20788 16528 20819
rect 17586 20816 17592 20828
rect 17644 20816 17650 20868
rect 17681 20859 17739 20865
rect 17681 20825 17693 20859
rect 17727 20856 17739 20859
rect 18785 20859 18843 20865
rect 18785 20856 18797 20859
rect 17727 20828 18797 20856
rect 17727 20825 17739 20828
rect 17681 20819 17739 20825
rect 18785 20825 18797 20828
rect 18831 20825 18843 20859
rect 18785 20819 18843 20825
rect 15160 20760 16528 20788
rect 15160 20748 15166 20760
rect 17494 20748 17500 20800
rect 17552 20788 17558 20800
rect 17865 20791 17923 20797
rect 17865 20788 17877 20791
rect 17552 20760 17877 20788
rect 17552 20748 17558 20760
rect 17865 20757 17877 20760
rect 17911 20788 17923 20791
rect 18322 20788 18328 20800
rect 17911 20760 18328 20788
rect 17911 20757 17923 20760
rect 17865 20751 17923 20757
rect 18322 20748 18328 20760
rect 18380 20748 18386 20800
rect 21450 20788 21456 20800
rect 21411 20760 21456 20788
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 21637 20791 21695 20797
rect 21637 20757 21649 20791
rect 21683 20788 21695 20791
rect 22922 20788 22928 20800
rect 21683 20760 22928 20788
rect 21683 20757 21695 20760
rect 21637 20751 21695 20757
rect 22922 20748 22928 20760
rect 22980 20748 22986 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 5902 20544 5908 20596
rect 5960 20584 5966 20596
rect 6454 20584 6460 20596
rect 5960 20556 6460 20584
rect 5960 20544 5966 20556
rect 6454 20544 6460 20556
rect 6512 20584 6518 20596
rect 6917 20587 6975 20593
rect 6917 20584 6929 20587
rect 6512 20556 6929 20584
rect 6512 20544 6518 20556
rect 6917 20553 6929 20556
rect 6963 20553 6975 20587
rect 6917 20547 6975 20553
rect 8570 20544 8576 20596
rect 8628 20584 8634 20596
rect 9582 20584 9588 20596
rect 8628 20556 9588 20584
rect 8628 20544 8634 20556
rect 9582 20544 9588 20556
rect 9640 20584 9646 20596
rect 9693 20587 9751 20593
rect 9693 20584 9705 20587
rect 9640 20556 9705 20584
rect 9640 20544 9646 20556
rect 9693 20553 9705 20556
rect 9739 20553 9751 20587
rect 9693 20547 9751 20553
rect 10689 20587 10747 20593
rect 10689 20553 10701 20587
rect 10735 20584 10747 20587
rect 10778 20584 10784 20596
rect 10735 20556 10784 20584
rect 10735 20553 10747 20556
rect 10689 20547 10747 20553
rect 10778 20544 10784 20556
rect 10836 20544 10842 20596
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11701 20587 11759 20593
rect 11701 20584 11713 20587
rect 11572 20556 11713 20584
rect 11572 20544 11578 20556
rect 11701 20553 11713 20556
rect 11747 20553 11759 20587
rect 11701 20547 11759 20553
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 13228 20556 14289 20584
rect 13228 20544 13234 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 15930 20584 15936 20596
rect 14792 20556 15936 20584
rect 14792 20544 14798 20556
rect 15930 20544 15936 20556
rect 15988 20584 15994 20596
rect 18690 20584 18696 20596
rect 15988 20556 18696 20584
rect 15988 20544 15994 20556
rect 18690 20544 18696 20556
rect 18748 20544 18754 20596
rect 20181 20587 20239 20593
rect 20181 20584 20193 20587
rect 19168 20556 20193 20584
rect 3050 20476 3056 20528
rect 3108 20516 3114 20528
rect 5442 20516 5448 20528
rect 3108 20488 5448 20516
rect 3108 20476 3114 20488
rect 2133 20451 2191 20457
rect 2133 20417 2145 20451
rect 2179 20448 2191 20451
rect 2222 20448 2228 20460
rect 2179 20420 2228 20448
rect 2179 20417 2191 20420
rect 2133 20411 2191 20417
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 2314 20408 2320 20460
rect 2372 20448 2378 20460
rect 3160 20457 3188 20488
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 5552 20488 7144 20516
rect 3145 20451 3203 20457
rect 2372 20420 2417 20448
rect 2372 20408 2378 20420
rect 3145 20417 3157 20451
rect 3191 20417 3203 20451
rect 3145 20411 3203 20417
rect 3878 20408 3884 20460
rect 3936 20448 3942 20460
rect 4065 20451 4123 20457
rect 4065 20448 4077 20451
rect 3936 20420 4077 20448
rect 3936 20408 3942 20420
rect 4065 20417 4077 20420
rect 4111 20417 4123 20451
rect 4246 20448 4252 20460
rect 4207 20420 4252 20448
rect 4065 20411 4123 20417
rect 4246 20408 4252 20420
rect 4304 20448 4310 20460
rect 4614 20448 4620 20460
rect 4304 20420 4620 20448
rect 4304 20408 4310 20420
rect 4614 20408 4620 20420
rect 4672 20408 4678 20460
rect 5258 20408 5264 20460
rect 5316 20448 5322 20460
rect 5552 20457 5580 20488
rect 5537 20451 5595 20457
rect 5537 20448 5549 20451
rect 5316 20420 5549 20448
rect 5316 20408 5322 20420
rect 5537 20417 5549 20420
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20448 6055 20451
rect 6086 20448 6092 20460
rect 6043 20420 6092 20448
rect 6043 20417 6055 20420
rect 5997 20411 6055 20417
rect 3418 20380 3424 20392
rect 3379 20352 3424 20380
rect 3418 20340 3424 20352
rect 3476 20340 3482 20392
rect 3970 20340 3976 20392
rect 4028 20380 4034 20392
rect 4341 20383 4399 20389
rect 4341 20380 4353 20383
rect 4028 20352 4353 20380
rect 4028 20340 4034 20352
rect 4341 20349 4353 20352
rect 4387 20349 4399 20383
rect 5828 20380 5856 20411
rect 6086 20408 6092 20420
rect 6144 20408 6150 20460
rect 7116 20457 7144 20488
rect 8478 20476 8484 20528
rect 8536 20516 8542 20528
rect 9493 20519 9551 20525
rect 9493 20516 9505 20519
rect 8536 20488 9505 20516
rect 8536 20476 8542 20488
rect 9493 20485 9505 20488
rect 9539 20485 9551 20519
rect 9493 20479 9551 20485
rect 11790 20476 11796 20528
rect 11848 20516 11854 20528
rect 15838 20516 15844 20528
rect 11848 20488 15844 20516
rect 11848 20476 11854 20488
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20417 7159 20451
rect 7374 20448 7380 20460
rect 7335 20420 7380 20448
rect 7101 20411 7159 20417
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20448 7619 20451
rect 8294 20448 8300 20460
rect 7607 20420 8300 20448
rect 7607 20417 7619 20420
rect 7561 20411 7619 20417
rect 8294 20408 8300 20420
rect 8352 20448 8358 20460
rect 9306 20448 9312 20460
rect 8352 20420 9312 20448
rect 8352 20408 8358 20420
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20448 10931 20451
rect 11054 20448 11060 20460
rect 10919 20420 11060 20448
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20448 11207 20451
rect 11698 20448 11704 20460
rect 11195 20420 11704 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20448 11943 20451
rect 11974 20448 11980 20460
rect 11931 20420 11980 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 12158 20448 12164 20460
rect 12119 20420 12164 20448
rect 12158 20408 12164 20420
rect 12216 20408 12222 20460
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 14274 20448 14280 20460
rect 12943 20420 14280 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 14274 20408 14280 20420
rect 14332 20408 14338 20460
rect 14568 20457 14596 20488
rect 15838 20476 15844 20488
rect 15896 20516 15902 20528
rect 19168 20516 19196 20556
rect 20181 20553 20193 20556
rect 20227 20584 20239 20587
rect 20809 20587 20867 20593
rect 20227 20556 20760 20584
rect 20227 20553 20239 20556
rect 20181 20547 20239 20553
rect 19981 20519 20039 20525
rect 19981 20516 19993 20519
rect 15896 20488 19196 20516
rect 15896 20476 15902 20488
rect 14553 20451 14611 20457
rect 14553 20417 14565 20451
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20448 14795 20451
rect 14826 20448 14832 20460
rect 14783 20420 14832 20448
rect 14783 20417 14795 20420
rect 14737 20411 14795 20417
rect 14826 20408 14832 20420
rect 14884 20408 14890 20460
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 15654 20448 15660 20460
rect 15611 20420 15660 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 15746 20408 15752 20460
rect 15804 20448 15810 20460
rect 15804 20420 15849 20448
rect 15804 20408 15810 20420
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 15988 20420 16033 20448
rect 15988 20408 15994 20420
rect 16298 20408 16304 20460
rect 16356 20448 16362 20460
rect 17770 20448 17776 20460
rect 16356 20420 16401 20448
rect 17731 20420 17776 20448
rect 16356 20408 16362 20420
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 19168 20457 19196 20488
rect 19306 20488 19993 20516
rect 19306 20460 19334 20488
rect 19981 20485 19993 20488
rect 20027 20516 20039 20519
rect 20732 20516 20760 20556
rect 20809 20553 20821 20587
rect 20855 20584 20867 20587
rect 21450 20584 21456 20596
rect 20855 20556 21456 20584
rect 20855 20553 20867 20556
rect 20809 20547 20867 20553
rect 21450 20544 21456 20556
rect 21508 20544 21514 20596
rect 20027 20488 20484 20516
rect 20732 20488 21312 20516
rect 20027 20485 20039 20488
rect 19981 20479 20039 20485
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 19153 20451 19211 20457
rect 19153 20417 19165 20451
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 6822 20380 6828 20392
rect 5828 20352 6828 20380
rect 4341 20343 4399 20349
rect 6104 20324 6132 20352
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7466 20340 7472 20392
rect 7524 20380 7530 20392
rect 10686 20380 10692 20392
rect 7524 20352 10692 20380
rect 7524 20340 7530 20352
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 11900 20352 12081 20380
rect 11900 20324 11928 20352
rect 12069 20349 12081 20352
rect 12115 20349 12127 20383
rect 12069 20343 12127 20349
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13170 20380 13176 20392
rect 13035 20352 13176 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 13170 20340 13176 20352
rect 13228 20340 13234 20392
rect 14458 20380 14464 20392
rect 14419 20352 14464 20380
rect 14458 20340 14464 20352
rect 14516 20340 14522 20392
rect 14642 20380 14648 20392
rect 14603 20352 14648 20380
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 18524 20380 18552 20411
rect 18064 20352 18552 20380
rect 18064 20324 18092 20352
rect 3050 20272 3056 20324
rect 3108 20312 3114 20324
rect 3329 20315 3387 20321
rect 3329 20312 3341 20315
rect 3108 20284 3341 20312
rect 3108 20272 3114 20284
rect 3329 20281 3341 20284
rect 3375 20281 3387 20315
rect 3329 20275 3387 20281
rect 6086 20272 6092 20324
rect 6144 20272 6150 20324
rect 9858 20312 9864 20324
rect 9771 20284 9864 20312
rect 9858 20272 9864 20284
rect 9916 20312 9922 20324
rect 10962 20312 10968 20324
rect 9916 20284 10968 20312
rect 9916 20272 9922 20284
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 11882 20272 11888 20324
rect 11940 20272 11946 20324
rect 11974 20272 11980 20324
rect 12032 20312 12038 20324
rect 12032 20284 12077 20312
rect 12032 20272 12038 20284
rect 14918 20272 14924 20324
rect 14976 20312 14982 20324
rect 16298 20312 16304 20324
rect 14976 20284 16304 20312
rect 14976 20272 14982 20284
rect 16298 20272 16304 20284
rect 16356 20312 16362 20324
rect 17957 20315 18015 20321
rect 17957 20312 17969 20315
rect 16356 20284 17969 20312
rect 16356 20272 16362 20284
rect 17957 20281 17969 20284
rect 18003 20312 18015 20315
rect 18046 20312 18052 20324
rect 18003 20284 18052 20312
rect 18003 20281 18015 20284
rect 17957 20275 18015 20281
rect 18046 20272 18052 20284
rect 18104 20272 18110 20324
rect 18138 20272 18144 20324
rect 18196 20312 18202 20324
rect 18708 20312 18736 20411
rect 19242 20408 19248 20460
rect 19300 20448 19334 20460
rect 19300 20420 19345 20448
rect 19300 20408 19306 20420
rect 18196 20284 18736 20312
rect 19352 20284 20208 20312
rect 18196 20272 18202 20284
rect 2130 20244 2136 20256
rect 2091 20216 2136 20244
rect 2130 20204 2136 20216
rect 2188 20204 2194 20256
rect 3234 20244 3240 20256
rect 3195 20216 3240 20244
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 3881 20247 3939 20253
rect 3881 20213 3893 20247
rect 3927 20244 3939 20247
rect 4062 20244 4068 20256
rect 3927 20216 4068 20244
rect 3927 20213 3939 20216
rect 3881 20207 3939 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5353 20247 5411 20253
rect 5353 20213 5365 20247
rect 5399 20244 5411 20247
rect 5626 20244 5632 20256
rect 5399 20216 5632 20244
rect 5399 20213 5411 20216
rect 5353 20207 5411 20213
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 9674 20244 9680 20256
rect 9635 20216 9680 20244
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 11054 20244 11060 20256
rect 11015 20216 11060 20244
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13265 20247 13323 20253
rect 13265 20244 13277 20247
rect 13136 20216 13277 20244
rect 13136 20204 13142 20216
rect 13265 20213 13277 20216
rect 13311 20213 13323 20247
rect 13265 20207 13323 20213
rect 14550 20204 14556 20256
rect 14608 20244 14614 20256
rect 15565 20247 15623 20253
rect 15565 20244 15577 20247
rect 14608 20216 15577 20244
rect 14608 20204 14614 20216
rect 15565 20213 15577 20216
rect 15611 20213 15623 20247
rect 15565 20207 15623 20213
rect 15654 20204 15660 20256
rect 15712 20244 15718 20256
rect 15838 20244 15844 20256
rect 15712 20216 15844 20244
rect 15712 20204 15718 20216
rect 15838 20204 15844 20216
rect 15896 20244 15902 20256
rect 17862 20244 17868 20256
rect 15896 20216 17868 20244
rect 15896 20204 15902 20216
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 18598 20244 18604 20256
rect 18559 20216 18604 20244
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 19352 20253 19380 20284
rect 20180 20256 20208 20284
rect 19337 20247 19395 20253
rect 19337 20213 19349 20247
rect 19383 20213 19395 20247
rect 19337 20207 19395 20213
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19521 20247 19579 20253
rect 19521 20244 19533 20247
rect 19484 20216 19533 20244
rect 19484 20204 19490 20216
rect 19521 20213 19533 20216
rect 19567 20213 19579 20247
rect 20162 20244 20168 20256
rect 20123 20216 20168 20244
rect 19521 20207 19579 20213
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20346 20244 20352 20256
rect 20307 20216 20352 20244
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 20456 20244 20484 20488
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 20990 20448 20996 20460
rect 20588 20420 20996 20448
rect 20588 20408 20594 20420
rect 20990 20408 20996 20420
rect 21048 20408 21054 20460
rect 21284 20457 21312 20488
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 21358 20448 21364 20460
rect 21315 20420 21364 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20417 22155 20451
rect 22922 20448 22928 20460
rect 22883 20420 22928 20448
rect 22097 20411 22155 20417
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 21085 20383 21143 20389
rect 21085 20380 21097 20383
rect 20956 20352 21097 20380
rect 20956 20340 20962 20352
rect 21085 20349 21097 20352
rect 21131 20349 21143 20383
rect 21085 20343 21143 20349
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20349 21235 20383
rect 21177 20343 21235 20349
rect 21192 20244 21220 20343
rect 21266 20272 21272 20324
rect 21324 20312 21330 20324
rect 22112 20312 22140 20411
rect 22922 20408 22928 20420
rect 22980 20408 22986 20460
rect 21324 20284 22140 20312
rect 21324 20272 21330 20284
rect 20456 20216 21220 20244
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 22189 20247 22247 20253
rect 22189 20244 22201 20247
rect 22152 20216 22201 20244
rect 22152 20204 22158 20216
rect 22189 20213 22201 20216
rect 22235 20213 22247 20247
rect 22738 20244 22744 20256
rect 22699 20216 22744 20244
rect 22189 20207 22247 20213
rect 22738 20204 22744 20216
rect 22796 20204 22802 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 2222 20000 2228 20052
rect 2280 20040 2286 20052
rect 3973 20043 4031 20049
rect 3973 20040 3985 20043
rect 2280 20012 3985 20040
rect 2280 20000 2286 20012
rect 3973 20009 3985 20012
rect 4019 20009 4031 20043
rect 3973 20003 4031 20009
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 4798 20040 4804 20052
rect 4571 20012 4804 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 4798 20000 4804 20012
rect 4856 20040 4862 20052
rect 5629 20043 5687 20049
rect 5629 20040 5641 20043
rect 4856 20012 5641 20040
rect 4856 20000 4862 20012
rect 5629 20009 5641 20012
rect 5675 20009 5687 20043
rect 5629 20003 5687 20009
rect 6270 20000 6276 20052
rect 6328 20040 6334 20052
rect 6365 20043 6423 20049
rect 6365 20040 6377 20043
rect 6328 20012 6377 20040
rect 6328 20000 6334 20012
rect 6365 20009 6377 20012
rect 6411 20009 6423 20043
rect 6365 20003 6423 20009
rect 6546 20000 6552 20052
rect 6604 20040 6610 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 6604 20012 6837 20040
rect 6604 20000 6610 20012
rect 6825 20009 6837 20012
rect 6871 20009 6883 20043
rect 6825 20003 6883 20009
rect 7374 20000 7380 20052
rect 7432 20040 7438 20052
rect 8297 20043 8355 20049
rect 8297 20040 8309 20043
rect 7432 20012 8309 20040
rect 7432 20000 7438 20012
rect 8297 20009 8309 20012
rect 8343 20009 8355 20043
rect 8297 20003 8355 20009
rect 2958 19972 2964 19984
rect 2919 19944 2964 19972
rect 2958 19932 2964 19944
rect 3016 19932 3022 19984
rect 3234 19864 3240 19916
rect 3292 19904 3298 19916
rect 6454 19904 6460 19916
rect 3292 19876 4660 19904
rect 6415 19876 6460 19904
rect 3292 19864 3298 19876
rect 1581 19839 1639 19845
rect 1581 19805 1593 19839
rect 1627 19805 1639 19839
rect 1581 19799 1639 19805
rect 1848 19839 1906 19845
rect 1848 19805 1860 19839
rect 1894 19836 1906 19839
rect 2130 19836 2136 19848
rect 1894 19808 2136 19836
rect 1894 19805 1906 19808
rect 1848 19799 1906 19805
rect 1596 19768 1624 19799
rect 2130 19796 2136 19808
rect 2188 19796 2194 19848
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 4632 19845 4660 19876
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 7650 19904 7656 19916
rect 7300 19876 7656 19904
rect 4098 19839 4156 19845
rect 4098 19836 4110 19839
rect 3476 19808 4110 19836
rect 3476 19796 3482 19808
rect 4098 19805 4110 19808
rect 4144 19805 4156 19839
rect 4098 19799 4156 19805
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 6362 19836 6368 19848
rect 4663 19808 5488 19836
rect 6323 19808 6368 19836
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 4890 19768 4896 19780
rect 1596 19740 4896 19768
rect 1872 19712 1900 19740
rect 4890 19728 4896 19740
rect 4948 19728 4954 19780
rect 1854 19660 1860 19712
rect 1912 19660 1918 19712
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 4157 19703 4215 19709
rect 4157 19700 4169 19703
rect 4120 19672 4169 19700
rect 4120 19660 4126 19672
rect 4157 19669 4169 19672
rect 4203 19669 4215 19703
rect 5460 19700 5488 19808
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 6546 19796 6552 19848
rect 6604 19836 6610 19848
rect 7300 19845 7328 19876
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 8312 19904 8340 20003
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11977 20043 12035 20049
rect 11977 20040 11989 20043
rect 11112 20012 11989 20040
rect 11112 20000 11118 20012
rect 11977 20009 11989 20012
rect 12023 20009 12035 20043
rect 11977 20003 12035 20009
rect 15746 20000 15752 20052
rect 15804 20040 15810 20052
rect 16117 20043 16175 20049
rect 16117 20040 16129 20043
rect 15804 20012 16129 20040
rect 15804 20000 15810 20012
rect 16117 20009 16129 20012
rect 16163 20009 16175 20043
rect 18138 20040 18144 20052
rect 16117 20003 16175 20009
rect 16316 20012 18144 20040
rect 8478 19972 8484 19984
rect 8439 19944 8484 19972
rect 8478 19932 8484 19944
rect 8536 19932 8542 19984
rect 10594 19932 10600 19984
rect 10652 19972 10658 19984
rect 11517 19975 11575 19981
rect 10652 19944 11468 19972
rect 10652 19932 10658 19944
rect 9401 19907 9459 19913
rect 9401 19904 9413 19907
rect 8312 19876 9413 19904
rect 9401 19873 9413 19876
rect 9447 19873 9459 19907
rect 9401 19867 9459 19873
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 11057 19907 11115 19913
rect 11057 19904 11069 19907
rect 9640 19876 11069 19904
rect 9640 19864 9646 19876
rect 11057 19873 11069 19876
rect 11103 19873 11115 19907
rect 11440 19904 11468 19944
rect 11517 19941 11529 19975
rect 11563 19972 11575 19975
rect 11882 19972 11888 19984
rect 11563 19944 11888 19972
rect 11563 19941 11575 19944
rect 11517 19935 11575 19941
rect 11882 19932 11888 19944
rect 11940 19932 11946 19984
rect 14918 19972 14924 19984
rect 12820 19944 14924 19972
rect 12820 19904 12848 19944
rect 14918 19932 14924 19944
rect 14976 19932 14982 19984
rect 14734 19904 14740 19916
rect 11440 19876 12848 19904
rect 12912 19876 14740 19904
rect 11057 19867 11115 19873
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 6604 19808 6653 19836
rect 6604 19796 6610 19808
rect 6641 19805 6653 19808
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7466 19836 7472 19848
rect 7427 19808 7472 19836
rect 7285 19799 7343 19805
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 7668 19836 7696 19864
rect 9125 19839 9183 19845
rect 7668 19808 8248 19836
rect 5537 19771 5595 19777
rect 5537 19737 5549 19771
rect 5583 19768 5595 19771
rect 5718 19768 5724 19780
rect 5583 19740 5724 19768
rect 5583 19737 5595 19740
rect 5537 19731 5595 19737
rect 5718 19728 5724 19740
rect 5776 19768 5782 19780
rect 7377 19771 7435 19777
rect 7377 19768 7389 19771
rect 5776 19740 7389 19768
rect 5776 19728 5782 19740
rect 7377 19737 7389 19740
rect 7423 19737 7435 19771
rect 7377 19731 7435 19737
rect 7742 19728 7748 19780
rect 7800 19768 7806 19780
rect 8113 19771 8171 19777
rect 8113 19768 8125 19771
rect 7800 19740 8125 19768
rect 7800 19728 7806 19740
rect 8113 19737 8125 19740
rect 8159 19737 8171 19771
rect 8220 19768 8248 19808
rect 9125 19805 9137 19839
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 11149 19839 11207 19845
rect 11149 19805 11161 19839
rect 11195 19836 11207 19839
rect 11790 19836 11796 19848
rect 11195 19808 11796 19836
rect 11195 19805 11207 19808
rect 11149 19799 11207 19805
rect 8313 19771 8371 19777
rect 8313 19768 8325 19771
rect 8220 19740 8325 19768
rect 8113 19731 8171 19737
rect 8313 19737 8325 19740
rect 8359 19737 8371 19771
rect 9140 19768 9168 19799
rect 11790 19796 11796 19808
rect 11848 19796 11854 19848
rect 11974 19836 11980 19848
rect 11935 19808 11980 19836
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 12124 19808 12173 19836
rect 12124 19796 12130 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 12912 19836 12940 19876
rect 14734 19864 14740 19876
rect 14792 19904 14798 19916
rect 15381 19907 15439 19913
rect 14792 19876 14872 19904
rect 14792 19864 14798 19876
rect 13078 19836 13084 19848
rect 12768 19808 12940 19836
rect 13039 19808 13084 19836
rect 12768 19796 12774 19808
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13262 19845 13268 19848
rect 13229 19839 13268 19845
rect 13229 19805 13241 19839
rect 13229 19799 13268 19805
rect 13262 19796 13268 19799
rect 13320 19796 13326 19848
rect 13587 19839 13645 19845
rect 13587 19805 13599 19839
rect 13633 19836 13645 19839
rect 13722 19836 13728 19848
rect 13633 19808 13728 19836
rect 13633 19805 13645 19808
rect 13587 19799 13645 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 9398 19768 9404 19780
rect 8313 19731 8371 19737
rect 8404 19740 8616 19768
rect 9140 19740 9404 19768
rect 8404 19700 8432 19740
rect 5460 19672 8432 19700
rect 8588 19700 8616 19740
rect 9398 19728 9404 19740
rect 9456 19728 9462 19780
rect 11992 19700 12020 19796
rect 13354 19768 13360 19780
rect 13315 19740 13360 19768
rect 13354 19728 13360 19740
rect 13412 19728 13418 19780
rect 13449 19771 13507 19777
rect 13449 19737 13461 19771
rect 13495 19768 13507 19771
rect 13814 19768 13820 19780
rect 13495 19740 13820 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 13814 19728 13820 19740
rect 13872 19768 13878 19780
rect 14844 19768 14872 19876
rect 15381 19873 15393 19907
rect 15427 19904 15439 19907
rect 15764 19904 15792 20000
rect 16316 19984 16344 20012
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 18322 20040 18328 20052
rect 18283 20012 18328 20040
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 20346 20040 20352 20052
rect 19935 20012 20352 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 21082 20000 21088 20052
rect 21140 20040 21146 20052
rect 21269 20043 21327 20049
rect 21269 20040 21281 20043
rect 21140 20012 21281 20040
rect 21140 20000 21146 20012
rect 21269 20009 21281 20012
rect 21315 20009 21327 20043
rect 21269 20003 21327 20009
rect 21358 20000 21364 20052
rect 21416 20040 21422 20052
rect 23385 20043 23443 20049
rect 23385 20040 23397 20043
rect 21416 20012 23397 20040
rect 21416 20000 21422 20012
rect 23385 20009 23397 20012
rect 23431 20009 23443 20043
rect 23385 20003 23443 20009
rect 16209 19975 16267 19981
rect 16209 19941 16221 19975
rect 16255 19972 16267 19975
rect 16298 19972 16304 19984
rect 16255 19944 16304 19972
rect 16255 19941 16267 19944
rect 16209 19935 16267 19941
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 20070 19972 20076 19984
rect 20031 19944 20076 19972
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 15427 19876 15792 19904
rect 15427 19873 15439 19876
rect 15381 19867 15439 19873
rect 15930 19864 15936 19916
rect 15988 19904 15994 19916
rect 16393 19907 16451 19913
rect 15988 19876 16160 19904
rect 15988 19864 15994 19876
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 15252 19808 15485 19836
rect 15252 19796 15258 19808
rect 15473 19805 15485 19808
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19836 15715 19839
rect 16022 19836 16028 19848
rect 15703 19808 16028 19836
rect 15703 19805 15715 19808
rect 15657 19799 15715 19805
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 16132 19845 16160 19876
rect 16393 19873 16405 19907
rect 16439 19904 16451 19907
rect 16758 19904 16764 19916
rect 16439 19876 16764 19904
rect 16439 19873 16451 19876
rect 16393 19867 16451 19873
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 16942 19904 16948 19916
rect 16903 19876 16948 19904
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 19705 19907 19763 19913
rect 19705 19904 19717 19907
rect 18656 19876 19717 19904
rect 18656 19864 18662 19876
rect 19705 19873 19717 19876
rect 19751 19873 19763 19907
rect 20364 19904 20392 20000
rect 20530 19904 20536 19916
rect 20364 19876 20536 19904
rect 19705 19867 19763 19873
rect 20530 19864 20536 19876
rect 20588 19904 20594 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20588 19876 20913 19904
rect 20588 19864 20594 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 19426 19836 19432 19848
rect 19387 19808 19432 19836
rect 16117 19799 16175 19805
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 14921 19771 14979 19777
rect 14921 19768 14933 19771
rect 13872 19740 14504 19768
rect 14844 19740 14933 19768
rect 13872 19728 13878 19740
rect 8588 19672 12020 19700
rect 13725 19703 13783 19709
rect 4157 19663 4215 19669
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 14274 19700 14280 19712
rect 13771 19672 14280 19700
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 14476 19700 14504 19740
rect 14921 19737 14933 19740
rect 14967 19737 14979 19771
rect 14921 19731 14979 19737
rect 17212 19771 17270 19777
rect 17212 19737 17224 19771
rect 17258 19768 17270 19771
rect 17678 19768 17684 19780
rect 17258 19740 17684 19768
rect 17258 19737 17270 19740
rect 17212 19731 17270 19737
rect 17678 19728 17684 19740
rect 17736 19728 17742 19780
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 17920 19740 19288 19768
rect 17920 19728 17926 19740
rect 16206 19700 16212 19712
rect 14476 19672 16212 19700
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 16298 19660 16304 19712
rect 16356 19700 16362 19712
rect 18414 19700 18420 19712
rect 16356 19672 18420 19700
rect 16356 19660 16362 19672
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 19260 19700 19288 19740
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 19904 19768 19932 19799
rect 20622 19796 20628 19848
rect 20680 19836 20686 19848
rect 20990 19836 20996 19848
rect 20680 19808 20996 19836
rect 20680 19796 20686 19808
rect 20990 19796 20996 19808
rect 21048 19836 21054 19848
rect 21085 19839 21143 19845
rect 21085 19836 21097 19839
rect 21048 19808 21097 19836
rect 21048 19796 21054 19808
rect 21085 19805 21097 19808
rect 21131 19805 21143 19839
rect 21085 19799 21143 19805
rect 21174 19796 21180 19848
rect 21232 19836 21238 19848
rect 22005 19839 22063 19845
rect 22005 19836 22017 19839
rect 21232 19808 22017 19836
rect 21232 19796 21238 19808
rect 22005 19805 22017 19808
rect 22051 19805 22063 19839
rect 22005 19799 22063 19805
rect 22272 19839 22330 19845
rect 22272 19805 22284 19839
rect 22318 19836 22330 19839
rect 22738 19836 22744 19848
rect 22318 19808 22744 19836
rect 22318 19805 22330 19808
rect 22272 19799 22330 19805
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 19392 19740 19932 19768
rect 19392 19728 19398 19740
rect 21266 19700 21272 19712
rect 19260 19672 21272 19700
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3513 19499 3571 19505
rect 3513 19465 3525 19499
rect 3559 19496 3571 19499
rect 3970 19496 3976 19508
rect 3559 19468 3976 19496
rect 3559 19465 3571 19468
rect 3513 19459 3571 19465
rect 3970 19456 3976 19468
rect 4028 19496 4034 19508
rect 5353 19499 5411 19505
rect 4028 19468 4384 19496
rect 4028 19456 4034 19468
rect 1673 19431 1731 19437
rect 1673 19397 1685 19431
rect 1719 19428 1731 19431
rect 1946 19428 1952 19440
rect 1719 19400 1952 19428
rect 1719 19397 1731 19400
rect 1673 19391 1731 19397
rect 1946 19388 1952 19400
rect 2004 19428 2010 19440
rect 4356 19437 4384 19468
rect 5353 19465 5365 19499
rect 5399 19496 5411 19499
rect 5442 19496 5448 19508
rect 5399 19468 5448 19496
rect 5399 19465 5411 19468
rect 5353 19459 5411 19465
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 8294 19496 8300 19508
rect 7484 19468 8300 19496
rect 4341 19431 4399 19437
rect 2004 19400 4292 19428
rect 2004 19388 2010 19400
rect 3142 19360 3148 19372
rect 3103 19332 3148 19360
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 4264 19360 4292 19400
rect 4341 19397 4353 19431
rect 4387 19397 4399 19431
rect 4341 19391 4399 19397
rect 4557 19431 4615 19437
rect 4557 19397 4569 19431
rect 4603 19428 4615 19431
rect 4706 19428 4712 19440
rect 4603 19400 4712 19428
rect 4603 19397 4615 19400
rect 4557 19391 4615 19397
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 5994 19428 6000 19440
rect 4816 19400 6000 19428
rect 4816 19360 4844 19400
rect 5994 19388 6000 19400
rect 6052 19388 6058 19440
rect 5258 19360 5264 19372
rect 4264 19332 4844 19360
rect 5219 19332 5264 19360
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 6546 19360 6552 19372
rect 5684 19332 6552 19360
rect 5684 19320 5690 19332
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 7484 19369 7512 19468
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 14826 19496 14832 19508
rect 13320 19468 13584 19496
rect 14787 19468 14832 19496
rect 13320 19456 13326 19468
rect 7558 19388 7564 19440
rect 7616 19428 7622 19440
rect 12710 19428 12716 19440
rect 7616 19400 8800 19428
rect 7616 19388 7622 19400
rect 8772 19369 8800 19400
rect 9508 19400 12716 19428
rect 9508 19369 9536 19400
rect 12710 19388 12716 19400
rect 12768 19388 12774 19440
rect 13556 19428 13584 19468
rect 14826 19456 14832 19468
rect 14884 19456 14890 19508
rect 15654 19496 15660 19508
rect 14936 19468 15660 19496
rect 14936 19428 14964 19468
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 15746 19456 15752 19508
rect 15804 19496 15810 19508
rect 16025 19499 16083 19505
rect 16025 19496 16037 19499
rect 15804 19468 16037 19496
rect 15804 19456 15810 19468
rect 16025 19465 16037 19468
rect 16071 19465 16083 19499
rect 16025 19459 16083 19465
rect 16114 19456 16120 19508
rect 16172 19496 16178 19508
rect 16301 19499 16359 19505
rect 16301 19496 16313 19499
rect 16172 19468 16313 19496
rect 16172 19456 16178 19468
rect 16301 19465 16313 19468
rect 16347 19465 16359 19499
rect 18046 19496 18052 19508
rect 18007 19468 18052 19496
rect 16301 19459 16359 19465
rect 13556 19400 14964 19428
rect 6733 19363 6791 19369
rect 6733 19360 6745 19363
rect 6696 19332 6745 19360
rect 6696 19320 6702 19332
rect 6733 19329 6745 19332
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19329 7527 19363
rect 8573 19363 8631 19369
rect 8573 19360 8585 19363
rect 7469 19323 7527 19329
rect 7576 19332 8585 19360
rect 2958 19252 2964 19304
rect 3016 19292 3022 19304
rect 3053 19295 3111 19301
rect 3053 19292 3065 19295
rect 3016 19264 3065 19292
rect 3016 19252 3022 19264
rect 3053 19261 3065 19264
rect 3099 19261 3111 19295
rect 3053 19255 3111 19261
rect 5442 19252 5448 19304
rect 5500 19292 5506 19304
rect 5500 19264 7052 19292
rect 5500 19252 5506 19264
rect 1854 19224 1860 19236
rect 1815 19196 1860 19224
rect 1854 19184 1860 19196
rect 1912 19184 1918 19236
rect 4709 19227 4767 19233
rect 4709 19193 4721 19227
rect 4755 19224 4767 19227
rect 5534 19224 5540 19236
rect 4755 19196 5540 19224
rect 4755 19193 4767 19196
rect 4709 19187 4767 19193
rect 5534 19184 5540 19196
rect 5592 19184 5598 19236
rect 4525 19159 4583 19165
rect 4525 19125 4537 19159
rect 4571 19156 4583 19159
rect 4614 19156 4620 19168
rect 4571 19128 4620 19156
rect 4571 19125 4583 19128
rect 4525 19119 4583 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 5552 19156 5580 19184
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 5552 19128 6561 19156
rect 6549 19125 6561 19128
rect 6595 19156 6607 19159
rect 6730 19156 6736 19168
rect 6595 19128 6736 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 6914 19156 6920 19168
rect 6875 19128 6920 19156
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7024 19156 7052 19264
rect 7282 19252 7288 19304
rect 7340 19292 7346 19304
rect 7576 19292 7604 19332
rect 8573 19329 8585 19332
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 10919 19332 11008 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 8846 19292 8852 19304
rect 7340 19264 7604 19292
rect 8807 19264 8852 19292
rect 7340 19252 7346 19264
rect 8846 19252 8852 19264
rect 8904 19252 8910 19304
rect 9398 19292 9404 19304
rect 9359 19264 9404 19292
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 10980 19292 11008 19332
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 12802 19360 12808 19372
rect 11112 19332 11157 19360
rect 12763 19332 12808 19360
rect 11112 19320 11118 19332
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 13262 19360 13268 19372
rect 13223 19332 13268 19360
rect 13262 19320 13268 19332
rect 13320 19320 13326 19372
rect 13446 19360 13452 19372
rect 13407 19332 13452 19360
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 13556 19369 13584 19400
rect 15838 19388 15844 19440
rect 15896 19428 15902 19440
rect 15896 19400 16160 19428
rect 15896 19388 15902 19400
rect 13541 19363 13599 19369
rect 13541 19329 13553 19363
rect 13587 19329 13599 19363
rect 13814 19360 13820 19372
rect 13775 19332 13820 19360
rect 13541 19323 13599 19329
rect 13814 19320 13820 19332
rect 13872 19320 13878 19372
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 16132 19369 16160 19400
rect 15013 19363 15071 19369
rect 15013 19360 15025 19363
rect 14516 19332 15025 19360
rect 14516 19320 14522 19332
rect 15013 19329 15025 19332
rect 15059 19360 15071 19363
rect 15697 19360 15792 19364
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15059 19336 15792 19360
rect 15059 19332 15725 19336
rect 15059 19329 15071 19332
rect 15013 19323 15071 19329
rect 11238 19292 11244 19304
rect 10980 19264 11244 19292
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 13722 19292 13728 19304
rect 13683 19264 13728 19292
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 15286 19292 15292 19304
rect 15247 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15764 19301 15792 19336
rect 15856 19332 15945 19360
rect 15749 19295 15807 19301
rect 15749 19261 15761 19295
rect 15795 19261 15807 19295
rect 15749 19255 15807 19261
rect 10870 19224 10876 19236
rect 10831 19196 10876 19224
rect 10870 19184 10876 19196
rect 10928 19184 10934 19236
rect 15197 19227 15255 19233
rect 15197 19193 15209 19227
rect 15243 19224 15255 19227
rect 15856 19224 15884 19332
rect 15933 19329 15945 19332
rect 15979 19360 15991 19363
rect 16117 19363 16175 19369
rect 15979 19332 16068 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 16040 19292 16068 19332
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16316 19360 16344 19459
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 18138 19456 18144 19508
rect 18196 19496 18202 19508
rect 20254 19496 20260 19508
rect 18196 19468 20260 19496
rect 18196 19456 18202 19468
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 20763 19468 22232 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 18969 19431 19027 19437
rect 18969 19397 18981 19431
rect 19015 19428 19027 19431
rect 20162 19428 20168 19440
rect 19015 19400 20168 19428
rect 19015 19397 19027 19400
rect 18969 19391 19027 19397
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 20272 19428 20300 19456
rect 20622 19437 20628 19440
rect 20349 19431 20407 19437
rect 20349 19428 20361 19431
rect 20272 19400 20361 19428
rect 20349 19397 20361 19400
rect 20395 19397 20407 19431
rect 20349 19391 20407 19397
rect 20565 19431 20628 19437
rect 20565 19397 20577 19431
rect 20611 19397 20628 19431
rect 20565 19391 20628 19397
rect 20622 19388 20628 19391
rect 20680 19388 20686 19440
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16316 19332 16865 19360
rect 16117 19323 16175 19329
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19360 17095 19363
rect 17770 19360 17776 19372
rect 17083 19332 17776 19360
rect 17083 19329 17095 19332
rect 17037 19323 17095 19329
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 18138 19320 18144 19372
rect 18196 19360 18202 19372
rect 18690 19360 18696 19372
rect 18196 19332 18241 19360
rect 18651 19332 18696 19360
rect 18196 19320 18202 19332
rect 18690 19320 18696 19332
rect 18748 19360 18754 19372
rect 19334 19360 19340 19372
rect 18748 19332 19340 19360
rect 18748 19320 18754 19332
rect 19334 19320 19340 19332
rect 19392 19360 19398 19372
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 19392 19332 19441 19360
rect 19392 19320 19398 19332
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19360 19671 19363
rect 19659 19350 20484 19360
rect 20732 19350 20760 19459
rect 21453 19431 21511 19437
rect 21453 19397 21465 19431
rect 21499 19397 21511 19431
rect 21453 19391 21511 19397
rect 19659 19332 20760 19350
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 17586 19292 17592 19304
rect 16040 19264 17592 19292
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 17681 19295 17739 19301
rect 17681 19261 17693 19295
rect 17727 19292 17739 19295
rect 17862 19292 17868 19304
rect 17727 19264 17868 19292
rect 17727 19261 17739 19264
rect 17681 19255 17739 19261
rect 15243 19196 15884 19224
rect 16853 19227 16911 19233
rect 15243 19193 15255 19196
rect 15197 19187 15255 19193
rect 16853 19193 16865 19227
rect 16899 19224 16911 19227
rect 17696 19224 17724 19255
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 18966 19292 18972 19304
rect 18927 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 16899 19196 17724 19224
rect 18785 19227 18843 19233
rect 16899 19193 16911 19196
rect 16853 19187 16911 19193
rect 18785 19193 18797 19227
rect 18831 19224 18843 19227
rect 19628 19224 19656 19323
rect 20456 19322 20760 19332
rect 20990 19320 20996 19372
rect 21048 19360 21054 19372
rect 21177 19363 21235 19369
rect 21177 19360 21189 19363
rect 21048 19332 21189 19360
rect 21048 19320 21054 19332
rect 21177 19329 21189 19332
rect 21223 19360 21235 19363
rect 21358 19360 21364 19372
rect 21223 19332 21364 19360
rect 21223 19329 21235 19332
rect 21177 19323 21235 19329
rect 21358 19320 21364 19332
rect 21416 19320 21422 19372
rect 21468 19360 21496 19391
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21468 19332 22017 19360
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22094 19320 22100 19372
rect 22152 19320 22158 19372
rect 22204 19369 22232 19468
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19329 22247 19363
rect 22189 19323 22247 19329
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21269 19295 21327 19301
rect 21269 19292 21281 19295
rect 21140 19264 21281 19292
rect 21140 19252 21146 19264
rect 21269 19261 21281 19264
rect 21315 19261 21327 19295
rect 21269 19255 21327 19261
rect 21453 19295 21511 19301
rect 21453 19261 21465 19295
rect 21499 19292 21511 19295
rect 22112 19292 22140 19320
rect 21499 19264 22140 19292
rect 21499 19261 21511 19264
rect 21453 19255 21511 19261
rect 21468 19224 21496 19255
rect 18831 19196 19656 19224
rect 19720 19196 21496 19224
rect 18831 19193 18843 19196
rect 18785 19187 18843 19193
rect 7561 19159 7619 19165
rect 7561 19156 7573 19159
rect 7024 19128 7573 19156
rect 7561 19125 7573 19128
rect 7607 19125 7619 19159
rect 7926 19156 7932 19168
rect 7887 19128 7932 19156
rect 7561 19119 7619 19125
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8386 19156 8392 19168
rect 8347 19128 8392 19156
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 9769 19159 9827 19165
rect 9769 19125 9781 19159
rect 9815 19156 9827 19159
rect 11146 19156 11152 19168
rect 9815 19128 11152 19156
rect 9815 19125 9827 19128
rect 9769 19119 9827 19125
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 12618 19156 12624 19168
rect 12579 19128 12624 19156
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 13630 19156 13636 19168
rect 13591 19128 13636 19156
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 17310 19156 17316 19168
rect 13964 19128 17316 19156
rect 13964 19116 13970 19128
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19156 17923 19159
rect 17954 19156 17960 19168
rect 17911 19128 17960 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 19720 19156 19748 19196
rect 19024 19128 19748 19156
rect 19797 19159 19855 19165
rect 19024 19116 19030 19128
rect 19797 19125 19809 19159
rect 19843 19156 19855 19159
rect 20346 19156 20352 19168
rect 19843 19128 20352 19156
rect 19843 19125 19855 19128
rect 19797 19119 19855 19125
rect 20346 19116 20352 19128
rect 20404 19116 20410 19168
rect 20530 19156 20536 19168
rect 20491 19128 20536 19156
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 22002 19156 22008 19168
rect 21963 19128 22008 19156
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 38286 19156 38292 19168
rect 38247 19128 38292 19156
rect 38286 19116 38292 19128
rect 38344 19116 38350 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 3292 18924 3341 18952
rect 3292 18912 3298 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 5626 18952 5632 18964
rect 5587 18924 5632 18952
rect 3329 18915 3387 18921
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 6914 18952 6920 18964
rect 6503 18924 6920 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8389 18955 8447 18961
rect 8389 18952 8401 18955
rect 8352 18924 8401 18952
rect 8352 18912 8358 18924
rect 8389 18921 8401 18924
rect 8435 18921 8447 18955
rect 8389 18915 8447 18921
rect 8573 18955 8631 18961
rect 8573 18921 8585 18955
rect 8619 18952 8631 18955
rect 8846 18952 8852 18964
rect 8619 18924 8852 18952
rect 8619 18921 8631 18924
rect 8573 18915 8631 18921
rect 8404 18884 8432 18915
rect 8846 18912 8852 18924
rect 8904 18912 8910 18964
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 13688 18924 14289 18952
rect 13688 18912 13694 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 14737 18955 14795 18961
rect 14737 18921 14749 18955
rect 14783 18952 14795 18955
rect 15470 18952 15476 18964
rect 14783 18924 15476 18952
rect 14783 18921 14795 18924
rect 14737 18915 14795 18921
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 16942 18952 16948 18964
rect 15580 18924 16948 18952
rect 9355 18887 9413 18893
rect 9355 18884 9367 18887
rect 8404 18856 9367 18884
rect 9355 18853 9367 18856
rect 9401 18853 9413 18887
rect 9355 18847 9413 18853
rect 11057 18887 11115 18893
rect 11057 18853 11069 18887
rect 11103 18884 11115 18887
rect 11238 18884 11244 18896
rect 11103 18856 11244 18884
rect 11103 18853 11115 18856
rect 11057 18847 11115 18853
rect 11238 18844 11244 18856
rect 11296 18844 11302 18896
rect 12434 18844 12440 18896
rect 12492 18884 12498 18896
rect 12713 18887 12771 18893
rect 12713 18884 12725 18887
rect 12492 18856 12725 18884
rect 12492 18844 12498 18856
rect 12713 18853 12725 18856
rect 12759 18884 12771 18887
rect 15580 18884 15608 18924
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 17678 18952 17684 18964
rect 17639 18924 17684 18952
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 18693 18955 18751 18961
rect 18693 18952 18705 18955
rect 17828 18924 18705 18952
rect 17828 18912 17834 18924
rect 18693 18921 18705 18924
rect 18739 18921 18751 18955
rect 18693 18915 18751 18921
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19613 18955 19671 18961
rect 19613 18952 19625 18955
rect 19392 18924 19625 18952
rect 19392 18912 19398 18924
rect 19613 18921 19625 18924
rect 19659 18921 19671 18955
rect 19613 18915 19671 18921
rect 21358 18912 21364 18964
rect 21416 18952 21422 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 21416 18924 22569 18952
rect 21416 18912 21422 18924
rect 22557 18921 22569 18924
rect 22603 18921 22615 18955
rect 22557 18915 22615 18921
rect 12759 18856 15608 18884
rect 16025 18887 16083 18893
rect 12759 18853 12771 18856
rect 12713 18847 12771 18853
rect 16025 18853 16037 18887
rect 16071 18884 16083 18887
rect 16298 18884 16304 18896
rect 16071 18856 16304 18884
rect 16071 18853 16083 18856
rect 16025 18847 16083 18853
rect 16298 18844 16304 18856
rect 16356 18884 16362 18896
rect 16574 18884 16580 18896
rect 16356 18856 16580 18884
rect 16356 18844 16362 18856
rect 16574 18844 16580 18856
rect 16632 18844 16638 18896
rect 18138 18844 18144 18896
rect 18196 18844 18202 18896
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 19300 18856 20576 18884
rect 19300 18844 19306 18856
rect 3050 18776 3056 18828
rect 3108 18816 3114 18828
rect 5813 18819 5871 18825
rect 3108 18788 4568 18816
rect 3108 18776 3114 18788
rect 2958 18708 2964 18760
rect 3016 18748 3022 18760
rect 3237 18751 3295 18757
rect 3237 18748 3249 18751
rect 3016 18720 3249 18748
rect 3016 18708 3022 18720
rect 3237 18717 3249 18720
rect 3283 18717 3295 18751
rect 4430 18748 4436 18760
rect 4391 18720 4436 18748
rect 3237 18711 3295 18717
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 4540 18757 4568 18788
rect 5813 18785 5825 18819
rect 5859 18816 5871 18819
rect 6638 18816 6644 18828
rect 5859 18788 6644 18816
rect 5859 18785 5871 18788
rect 5813 18779 5871 18785
rect 6638 18776 6644 18788
rect 6696 18776 6702 18828
rect 7466 18816 7472 18828
rect 7379 18788 7472 18816
rect 7466 18776 7472 18788
rect 7524 18816 7530 18828
rect 7926 18816 7932 18828
rect 7524 18788 7932 18816
rect 7524 18776 7530 18788
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 10597 18819 10655 18825
rect 10597 18816 10609 18819
rect 9140 18788 10609 18816
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18717 4583 18751
rect 5534 18748 5540 18760
rect 5495 18720 5540 18748
rect 4525 18711 4583 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 7561 18751 7619 18757
rect 7561 18748 7573 18751
rect 6488 18720 7573 18748
rect 5902 18640 5908 18692
rect 5960 18680 5966 18692
rect 6273 18683 6331 18689
rect 6273 18680 6285 18683
rect 5960 18652 6285 18680
rect 5960 18640 5966 18652
rect 6273 18649 6285 18652
rect 6319 18649 6331 18683
rect 6273 18643 6331 18649
rect 4614 18572 4620 18624
rect 4672 18612 4678 18624
rect 6488 18621 6516 18720
rect 7561 18717 7573 18720
rect 7607 18748 7619 18751
rect 7650 18748 7656 18760
rect 7607 18720 7656 18748
rect 7607 18717 7619 18720
rect 7561 18711 7619 18717
rect 7650 18708 7656 18720
rect 7708 18708 7714 18760
rect 7742 18708 7748 18760
rect 7800 18708 7806 18760
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 9140 18757 9168 18788
rect 10597 18785 10609 18788
rect 10643 18785 10655 18819
rect 15286 18816 15292 18828
rect 10597 18779 10655 18785
rect 12406 18788 15292 18816
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 8168 18720 9137 18748
rect 8168 18708 8174 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18748 10747 18751
rect 12406 18748 12434 18788
rect 15286 18776 15292 18788
rect 15344 18816 15350 18828
rect 16390 18816 16396 18828
rect 15344 18788 16396 18816
rect 15344 18776 15350 18788
rect 16390 18776 16396 18788
rect 16448 18776 16454 18828
rect 18049 18819 18107 18825
rect 18049 18785 18061 18819
rect 18095 18816 18107 18819
rect 18156 18816 18184 18844
rect 18095 18788 20392 18816
rect 18095 18785 18107 18788
rect 18049 18779 18107 18785
rect 20364 18760 20392 18788
rect 10735 18720 12434 18748
rect 12529 18751 12587 18757
rect 10735 18717 10747 18720
rect 10689 18711 10747 18717
rect 12529 18717 12541 18751
rect 12575 18748 12587 18751
rect 12894 18748 12900 18760
rect 12575 18720 12900 18748
rect 12575 18717 12587 18720
rect 12529 18711 12587 18717
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 14090 18708 14096 18760
rect 14148 18748 14154 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 14148 18720 14473 18748
rect 14148 18708 14154 18720
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 15841 18751 15899 18757
rect 14608 18720 14653 18748
rect 14608 18708 14614 18720
rect 15841 18717 15853 18751
rect 15887 18748 15899 18751
rect 17770 18748 17776 18760
rect 15887 18720 17776 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18748 17923 18751
rect 17954 18748 17960 18760
rect 17911 18720 17960 18748
rect 17911 18717 17923 18720
rect 17865 18711 17923 18717
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 18138 18748 18144 18760
rect 18099 18720 18144 18748
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18598 18748 18604 18760
rect 18559 18720 18604 18748
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 20162 18748 20168 18760
rect 20123 18720 20168 18748
rect 20162 18708 20168 18720
rect 20220 18708 20226 18760
rect 20346 18748 20352 18760
rect 20307 18720 20352 18748
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 20548 18748 20576 18856
rect 21174 18748 21180 18760
rect 20548 18720 21180 18748
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 21444 18751 21502 18757
rect 21444 18717 21456 18751
rect 21490 18748 21502 18751
rect 22002 18748 22008 18760
rect 21490 18720 22008 18748
rect 21490 18717 21502 18720
rect 21444 18711 21502 18717
rect 22002 18708 22008 18720
rect 22060 18708 22066 18760
rect 7760 18680 7788 18708
rect 8205 18683 8263 18689
rect 8205 18680 8217 18683
rect 6656 18652 7604 18680
rect 7760 18652 8217 18680
rect 6656 18621 6684 18652
rect 7576 18624 7604 18652
rect 8205 18649 8217 18652
rect 8251 18680 8263 18683
rect 10778 18680 10784 18692
rect 8251 18652 10784 18680
rect 8251 18649 8263 18652
rect 8205 18643 8263 18649
rect 10778 18640 10784 18652
rect 10836 18640 10842 18692
rect 13357 18683 13415 18689
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 13630 18680 13636 18692
rect 13403 18652 13636 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13630 18640 13636 18652
rect 13688 18640 13694 18692
rect 13998 18680 14004 18692
rect 13832 18652 14004 18680
rect 4709 18615 4767 18621
rect 4709 18612 4721 18615
rect 4672 18584 4721 18612
rect 4672 18572 4678 18584
rect 4709 18581 4721 18584
rect 4755 18581 4767 18615
rect 4709 18575 4767 18581
rect 5813 18615 5871 18621
rect 5813 18581 5825 18615
rect 5859 18612 5871 18615
rect 6473 18615 6531 18621
rect 6473 18612 6485 18615
rect 5859 18584 6485 18612
rect 5859 18581 5871 18584
rect 5813 18575 5871 18581
rect 6473 18581 6485 18584
rect 6519 18581 6531 18615
rect 6473 18575 6531 18581
rect 6641 18615 6699 18621
rect 6641 18581 6653 18615
rect 6687 18581 6699 18615
rect 7098 18612 7104 18624
rect 7059 18584 7104 18612
rect 6641 18575 6699 18581
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 7558 18572 7564 18624
rect 7616 18572 7622 18624
rect 7745 18615 7803 18621
rect 7745 18581 7757 18615
rect 7791 18612 7803 18615
rect 7834 18612 7840 18624
rect 7791 18584 7840 18612
rect 7791 18581 7803 18584
rect 7745 18575 7803 18581
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 8415 18615 8473 18621
rect 8415 18581 8427 18615
rect 8461 18612 8473 18615
rect 9950 18612 9956 18624
rect 8461 18584 9956 18612
rect 8461 18581 8473 18584
rect 8415 18575 8473 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 13449 18615 13507 18621
rect 13449 18612 13461 18615
rect 12216 18584 13461 18612
rect 12216 18572 12222 18584
rect 13449 18581 13461 18584
rect 13495 18612 13507 18615
rect 13832 18612 13860 18652
rect 13998 18640 14004 18652
rect 14056 18640 14062 18692
rect 14274 18680 14280 18692
rect 14235 18652 14280 18680
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 17037 18683 17095 18689
rect 17037 18649 17049 18683
rect 17083 18680 17095 18683
rect 17494 18680 17500 18692
rect 17083 18652 17500 18680
rect 17083 18649 17095 18652
rect 17037 18643 17095 18649
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 17586 18640 17592 18692
rect 17644 18680 17650 18692
rect 19521 18683 19579 18689
rect 19521 18680 19533 18683
rect 17644 18652 19533 18680
rect 17644 18640 17650 18652
rect 19521 18649 19533 18652
rect 19567 18680 19579 18683
rect 20714 18680 20720 18692
rect 19567 18652 20720 18680
rect 19567 18649 19579 18652
rect 19521 18643 19579 18649
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 13495 18584 13860 18612
rect 13495 18581 13507 18584
rect 13449 18575 13507 18581
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 16482 18612 16488 18624
rect 13964 18584 16488 18612
rect 13964 18572 13970 18584
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 17126 18612 17132 18624
rect 17087 18584 17132 18612
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 20254 18612 20260 18624
rect 20215 18584 20260 18612
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 3881 18411 3939 18417
rect 3881 18377 3893 18411
rect 3927 18408 3939 18411
rect 4706 18408 4712 18420
rect 3927 18380 4712 18408
rect 3927 18377 3939 18380
rect 3881 18371 3939 18377
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 6917 18411 6975 18417
rect 6917 18408 6929 18411
rect 6328 18380 6929 18408
rect 6328 18368 6334 18380
rect 6917 18377 6929 18380
rect 6963 18377 6975 18411
rect 6917 18371 6975 18377
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 10137 18411 10195 18417
rect 10137 18408 10149 18411
rect 8168 18380 10149 18408
rect 8168 18368 8174 18380
rect 10137 18377 10149 18380
rect 10183 18377 10195 18411
rect 10778 18408 10784 18420
rect 10739 18380 10784 18408
rect 10137 18371 10195 18377
rect 10778 18368 10784 18380
rect 10836 18408 10842 18420
rect 13906 18408 13912 18420
rect 10836 18380 12434 18408
rect 10836 18368 10842 18380
rect 3237 18343 3295 18349
rect 3237 18309 3249 18343
rect 3283 18340 3295 18343
rect 5721 18343 5779 18349
rect 5721 18340 5733 18343
rect 3283 18312 4752 18340
rect 3283 18309 3295 18312
rect 3237 18303 3295 18309
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18272 3019 18275
rect 3881 18275 3939 18281
rect 3881 18272 3893 18275
rect 3007 18244 3893 18272
rect 3007 18241 3019 18244
rect 2961 18235 3019 18241
rect 3881 18241 3893 18244
rect 3927 18272 3939 18275
rect 4430 18272 4436 18284
rect 3927 18244 4436 18272
rect 3927 18241 3939 18244
rect 3881 18235 3939 18241
rect 4430 18232 4436 18244
rect 4488 18232 4494 18284
rect 4614 18272 4620 18284
rect 4575 18244 4620 18272
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 4724 18281 4752 18312
rect 5000 18312 5733 18340
rect 5000 18281 5028 18312
rect 5721 18309 5733 18312
rect 5767 18340 5779 18343
rect 6086 18340 6092 18352
rect 5767 18312 6092 18340
rect 5767 18309 5779 18312
rect 5721 18303 5779 18309
rect 6086 18300 6092 18312
rect 6144 18300 6150 18352
rect 6549 18343 6607 18349
rect 6549 18309 6561 18343
rect 6595 18340 6607 18343
rect 6638 18340 6644 18352
rect 6595 18312 6644 18340
rect 6595 18309 6607 18312
rect 6549 18303 6607 18309
rect 6638 18300 6644 18312
rect 6696 18300 6702 18352
rect 6765 18343 6823 18349
rect 6765 18309 6777 18343
rect 6811 18340 6823 18343
rect 7098 18340 7104 18352
rect 6811 18312 7104 18340
rect 6811 18309 6823 18312
rect 6765 18303 6823 18309
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 8386 18300 8392 18352
rect 8444 18340 8450 18352
rect 9002 18343 9060 18349
rect 9002 18340 9014 18343
rect 8444 18312 9014 18340
rect 8444 18300 8450 18312
rect 9002 18309 9014 18312
rect 9048 18309 9060 18343
rect 10686 18340 10692 18352
rect 10647 18312 10692 18340
rect 9002 18303 9060 18309
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 12406 18340 12434 18380
rect 13096 18380 13912 18408
rect 12805 18343 12863 18349
rect 12805 18340 12817 18343
rect 12406 18312 12817 18340
rect 12805 18309 12817 18312
rect 12851 18340 12863 18343
rect 12986 18340 12992 18352
rect 12851 18312 12992 18340
rect 12851 18309 12863 18312
rect 12805 18303 12863 18309
rect 12986 18300 12992 18312
rect 13044 18300 13050 18352
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 5534 18272 5540 18284
rect 5495 18244 5540 18272
rect 4985 18235 5043 18241
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8018 18272 8024 18284
rect 7979 18244 8024 18272
rect 8018 18232 8024 18244
rect 8076 18232 8082 18284
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 8478 18272 8484 18284
rect 8159 18244 8484 18272
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 11882 18272 11888 18284
rect 11843 18244 11888 18272
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 12621 18275 12679 18281
rect 12621 18272 12633 18275
rect 12124 18244 12633 18272
rect 12124 18232 12130 18244
rect 12621 18241 12633 18244
rect 12667 18272 12679 18275
rect 12710 18272 12716 18284
rect 12667 18244 12716 18272
rect 12667 18241 12679 18244
rect 12621 18235 12679 18241
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 3050 18204 3056 18216
rect 3011 18176 3056 18204
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 3237 18207 3295 18213
rect 3237 18173 3249 18207
rect 3283 18173 3295 18207
rect 3237 18167 3295 18173
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 5718 18204 5724 18216
rect 4939 18176 5724 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 3252 18136 3280 18167
rect 5718 18164 5724 18176
rect 5776 18164 5782 18216
rect 7926 18204 7932 18216
rect 7887 18176 7932 18204
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8757 18207 8815 18213
rect 8757 18204 8769 18207
rect 8260 18176 8769 18204
rect 8260 18164 8266 18176
rect 8757 18173 8769 18176
rect 8803 18173 8815 18207
rect 12158 18204 12164 18216
rect 12119 18176 12164 18204
rect 8757 18167 8815 18173
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 3878 18136 3884 18148
rect 3252 18108 3884 18136
rect 3878 18096 3884 18108
rect 3936 18136 3942 18148
rect 13096 18136 13124 18380
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 14090 18408 14096 18420
rect 14051 18380 14096 18408
rect 14090 18368 14096 18380
rect 14148 18368 14154 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 18417 18411 18475 18417
rect 18417 18408 18429 18411
rect 18380 18380 18429 18408
rect 18380 18368 18386 18380
rect 18417 18377 18429 18380
rect 18463 18408 18475 18411
rect 20438 18408 20444 18420
rect 18463 18380 20444 18408
rect 18463 18377 18475 18380
rect 18417 18371 18475 18377
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 15562 18300 15568 18352
rect 15620 18300 15626 18352
rect 17770 18340 17776 18352
rect 17683 18312 17776 18340
rect 17770 18300 17776 18312
rect 17828 18340 17834 18352
rect 19058 18340 19064 18352
rect 17828 18312 19064 18340
rect 17828 18300 17834 18312
rect 19058 18300 19064 18312
rect 19116 18300 19122 18352
rect 19604 18343 19662 18349
rect 19604 18309 19616 18343
rect 19650 18340 19662 18343
rect 20254 18340 20260 18352
rect 19650 18312 20260 18340
rect 19650 18309 19662 18312
rect 19604 18303 19662 18309
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 13464 18204 13492 18235
rect 13538 18232 13544 18284
rect 13596 18272 13602 18284
rect 13725 18275 13783 18281
rect 13596 18244 13641 18272
rect 13596 18232 13602 18244
rect 13725 18241 13737 18275
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 13740 18204 13768 18235
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 13998 18281 14004 18284
rect 13955 18275 14004 18281
rect 13872 18244 13917 18272
rect 13872 18232 13878 18244
rect 13955 18241 13967 18275
rect 14001 18241 14004 18275
rect 13955 18235 14004 18241
rect 13998 18232 14004 18235
rect 14056 18232 14062 18284
rect 15194 18272 15200 18284
rect 15155 18244 15200 18272
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15580 18272 15608 18300
rect 15304 18244 15608 18272
rect 15304 18216 15332 18244
rect 17494 18232 17500 18284
rect 17552 18272 17558 18284
rect 17589 18275 17647 18281
rect 17589 18272 17601 18275
rect 17552 18244 17601 18272
rect 17552 18232 17558 18244
rect 17589 18241 17601 18244
rect 17635 18272 17647 18275
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 17635 18244 18337 18272
rect 17635 18241 17647 18244
rect 17589 18235 17647 18241
rect 18325 18241 18337 18244
rect 18371 18272 18383 18275
rect 18598 18272 18604 18284
rect 18371 18244 18604 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 19337 18275 19395 18281
rect 19337 18241 19349 18275
rect 19383 18272 19395 18275
rect 19978 18272 19984 18284
rect 19383 18244 19984 18272
rect 19383 18241 19395 18244
rect 19337 18235 19395 18241
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 14090 18204 14096 18216
rect 13464 18176 13676 18204
rect 13740 18176 14096 18204
rect 3936 18108 7972 18136
rect 3936 18096 3942 18108
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 4798 18068 4804 18080
rect 4479 18040 4804 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 6730 18068 6736 18080
rect 6691 18040 6736 18068
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18068 7711 18071
rect 7834 18068 7840 18080
rect 7699 18040 7840 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 7944 18068 7972 18108
rect 9692 18108 13124 18136
rect 13648 18136 13676 18176
rect 14090 18164 14096 18176
rect 14148 18164 14154 18216
rect 15286 18204 15292 18216
rect 15199 18176 15292 18204
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 15565 18207 15623 18213
rect 15565 18204 15577 18207
rect 15436 18176 15577 18204
rect 15436 18164 15442 18176
rect 15565 18173 15577 18176
rect 15611 18173 15623 18207
rect 15565 18167 15623 18173
rect 17954 18136 17960 18148
rect 13648 18108 17960 18136
rect 9692 18068 9720 18108
rect 17954 18096 17960 18108
rect 18012 18096 18018 18148
rect 11698 18068 11704 18080
rect 7944 18040 9720 18068
rect 11659 18040 11704 18068
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 12986 18068 12992 18080
rect 12584 18040 12992 18068
rect 12584 18028 12590 18040
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 4614 17864 4620 17876
rect 4571 17836 4620 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 7745 17867 7803 17873
rect 7745 17833 7757 17867
rect 7791 17864 7803 17867
rect 7926 17864 7932 17876
rect 7791 17836 7932 17864
rect 7791 17833 7803 17836
rect 7745 17827 7803 17833
rect 7926 17824 7932 17836
rect 7984 17824 7990 17876
rect 12437 17867 12495 17873
rect 12437 17833 12449 17867
rect 12483 17864 12495 17867
rect 12526 17864 12532 17876
rect 12483 17836 12532 17864
rect 12483 17833 12495 17836
rect 12437 17827 12495 17833
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12621 17867 12679 17873
rect 12621 17833 12633 17867
rect 12667 17864 12679 17867
rect 12802 17864 12808 17876
rect 12667 17836 12808 17864
rect 12667 17833 12679 17836
rect 12621 17827 12679 17833
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 13081 17867 13139 17873
rect 13081 17833 13093 17867
rect 13127 17864 13139 17867
rect 13262 17864 13268 17876
rect 13127 17836 13268 17864
rect 13127 17833 13139 17836
rect 13081 17827 13139 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 13722 17864 13728 17876
rect 13372 17836 13728 17864
rect 6457 17799 6515 17805
rect 6457 17765 6469 17799
rect 6503 17796 6515 17799
rect 6638 17796 6644 17808
rect 6503 17768 6644 17796
rect 6503 17765 6515 17768
rect 6457 17759 6515 17765
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 10686 17756 10692 17808
rect 10744 17756 10750 17808
rect 13372 17796 13400 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15470 17824 15476 17876
rect 15528 17864 15534 17876
rect 17770 17864 17776 17876
rect 15528 17836 17776 17864
rect 15528 17824 15534 17836
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 17954 17864 17960 17876
rect 17915 17836 17960 17864
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 18138 17824 18144 17876
rect 18196 17864 18202 17876
rect 18601 17867 18659 17873
rect 18601 17864 18613 17867
rect 18196 17836 18613 17864
rect 18196 17824 18202 17836
rect 18601 17833 18613 17836
rect 18647 17833 18659 17867
rect 18601 17827 18659 17833
rect 11532 17768 13400 17796
rect 13541 17799 13599 17805
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 5534 17728 5540 17740
rect 4295 17700 5540 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 6181 17731 6239 17737
rect 6181 17697 6193 17731
rect 6227 17728 6239 17731
rect 8110 17728 8116 17740
rect 6227 17700 8116 17728
rect 6227 17697 6239 17700
rect 6181 17691 6239 17697
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10704 17728 10732 17756
rect 11532 17740 11560 17768
rect 13541 17765 13553 17799
rect 13587 17796 13599 17799
rect 13630 17796 13636 17808
rect 13587 17768 13636 17796
rect 13587 17765 13599 17768
rect 13541 17759 13599 17765
rect 13630 17756 13636 17768
rect 13688 17756 13694 17808
rect 14458 17756 14464 17808
rect 14516 17796 14522 17808
rect 15841 17799 15899 17805
rect 15841 17796 15853 17799
rect 14516 17768 15853 17796
rect 14516 17756 14522 17768
rect 15841 17765 15853 17768
rect 15887 17765 15899 17799
rect 18230 17796 18236 17808
rect 15841 17759 15899 17765
rect 17604 17768 18236 17796
rect 11514 17728 11520 17740
rect 10091 17700 10732 17728
rect 11427 17700 11520 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 14090 17728 14096 17740
rect 13280 17700 14096 17728
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 4157 17663 4215 17669
rect 4157 17660 4169 17663
rect 3283 17632 4169 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 4157 17629 4169 17632
rect 4203 17660 4215 17663
rect 4706 17660 4712 17672
rect 4203 17632 4712 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 4985 17663 5043 17669
rect 4985 17660 4997 17663
rect 4856 17632 4997 17660
rect 4856 17620 4862 17632
rect 4985 17629 4997 17632
rect 5031 17629 5043 17663
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 4985 17623 5043 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5258 17620 5264 17672
rect 5316 17660 5322 17672
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 5316 17632 6101 17660
rect 5316 17620 5322 17632
rect 6089 17629 6101 17632
rect 6135 17660 6147 17663
rect 6730 17660 6736 17672
rect 6135 17632 6736 17660
rect 6135 17629 6147 17632
rect 6089 17623 6147 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 7098 17620 7104 17672
rect 7156 17660 7162 17672
rect 7341 17663 7399 17669
rect 7341 17660 7353 17663
rect 7156 17632 7353 17660
rect 7156 17620 7162 17632
rect 7341 17629 7353 17632
rect 7387 17629 7399 17663
rect 7341 17623 7399 17629
rect 7459 17657 7517 17663
rect 7459 17623 7471 17657
rect 7505 17623 7517 17657
rect 3142 17552 3148 17604
rect 3200 17592 3206 17604
rect 3421 17595 3479 17601
rect 3421 17592 3433 17595
rect 3200 17564 3433 17592
rect 3200 17552 3206 17564
rect 3421 17561 3433 17564
rect 3467 17592 3479 17595
rect 5276 17592 5304 17620
rect 7459 17617 7517 17623
rect 7561 17660 7619 17663
rect 7650 17660 7656 17672
rect 7561 17657 7656 17660
rect 7561 17623 7573 17657
rect 7607 17632 7656 17657
rect 7607 17623 7619 17632
rect 7561 17617 7619 17623
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17660 10287 17663
rect 10594 17660 10600 17672
rect 10275 17632 10600 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 12066 17660 12072 17672
rect 11287 17632 12072 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 13170 17620 13176 17672
rect 13228 17660 13234 17672
rect 13280 17669 13308 17700
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 15151 17700 16221 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 16209 17697 16221 17700
rect 16255 17728 16267 17731
rect 16850 17728 16856 17740
rect 16255 17700 16856 17728
rect 16255 17697 16267 17700
rect 16209 17691 16267 17697
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 13265 17663 13323 17669
rect 13265 17660 13277 17663
rect 13228 17632 13277 17660
rect 13228 17620 13234 17632
rect 13265 17629 13277 17632
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 13538 17660 13544 17672
rect 13403 17632 13544 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 13633 17663 13691 17669
rect 13633 17629 13645 17663
rect 13679 17660 13691 17663
rect 13814 17660 13820 17672
rect 13679 17632 13820 17660
rect 13679 17629 13691 17632
rect 13633 17623 13691 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 15010 17660 15016 17672
rect 14971 17632 15016 17660
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 16025 17663 16083 17669
rect 16025 17660 16037 17663
rect 15344 17632 16037 17660
rect 15344 17620 15350 17632
rect 16025 17629 16037 17632
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 16114 17620 16120 17672
rect 16172 17660 16178 17672
rect 16172 17632 16217 17660
rect 16172 17620 16178 17632
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 17604 17669 17632 17768
rect 18230 17756 18236 17768
rect 18288 17756 18294 17808
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 17589 17663 17647 17669
rect 16356 17632 16401 17660
rect 16356 17620 16362 17632
rect 17589 17629 17601 17663
rect 17635 17629 17647 17663
rect 17696 17660 17724 17691
rect 17696 17632 18460 17660
rect 17589 17623 17647 17629
rect 3467 17564 5304 17592
rect 3467 17561 3479 17564
rect 3421 17555 3479 17561
rect 7474 17536 7502 17617
rect 18432 17604 18460 17632
rect 11333 17595 11391 17601
rect 11333 17592 11345 17595
rect 10428 17564 11345 17592
rect 10428 17536 10456 17564
rect 11333 17561 11345 17564
rect 11379 17561 11391 17595
rect 11333 17555 11391 17561
rect 12253 17595 12311 17601
rect 12253 17561 12265 17595
rect 12299 17592 12311 17595
rect 15470 17592 15476 17604
rect 12299 17564 15476 17592
rect 12299 17561 12311 17564
rect 12253 17555 12311 17561
rect 15470 17552 15476 17564
rect 15528 17552 15534 17604
rect 18414 17592 18420 17604
rect 15672 17564 15976 17592
rect 18375 17564 18420 17592
rect 15672 17536 15700 17564
rect 5350 17524 5356 17536
rect 5311 17496 5356 17524
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 7466 17484 7472 17536
rect 7524 17484 7530 17536
rect 10410 17524 10416 17536
rect 10371 17496 10416 17524
rect 10410 17484 10416 17496
rect 10468 17484 10474 17536
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 10873 17527 10931 17533
rect 10873 17524 10885 17527
rect 10560 17496 10885 17524
rect 10560 17484 10566 17496
rect 10873 17493 10885 17496
rect 10919 17493 10931 17527
rect 10873 17487 10931 17493
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12453 17527 12511 17533
rect 12453 17524 12465 17527
rect 11756 17496 12465 17524
rect 11756 17484 11762 17496
rect 12453 17493 12465 17496
rect 12499 17493 12511 17527
rect 12453 17487 12511 17493
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 15654 17524 15660 17536
rect 13044 17496 15660 17524
rect 13044 17484 13050 17496
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 15948 17524 15976 17564
rect 18414 17552 18420 17564
rect 18472 17552 18478 17604
rect 18617 17527 18675 17533
rect 18617 17524 18629 17527
rect 15948 17496 18629 17524
rect 18617 17493 18629 17496
rect 18663 17493 18675 17527
rect 18782 17524 18788 17536
rect 18743 17496 18788 17524
rect 18617 17487 18675 17493
rect 18782 17484 18788 17496
rect 18840 17484 18846 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 4801 17323 4859 17329
rect 4801 17289 4813 17323
rect 4847 17320 4859 17323
rect 5534 17320 5540 17332
rect 4847 17292 5540 17320
rect 4847 17289 4859 17292
rect 4801 17283 4859 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 7098 17320 7104 17332
rect 7059 17292 7104 17320
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 9824 17292 10640 17320
rect 9824 17280 9830 17292
rect 3436 17224 5120 17252
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 3436 17125 3464 17224
rect 3688 17187 3746 17193
rect 3688 17153 3700 17187
rect 3734 17184 3746 17187
rect 4062 17184 4068 17196
rect 3734 17156 4068 17184
rect 3734 17153 3746 17156
rect 3688 17147 3746 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 5092 17184 5120 17224
rect 5166 17212 5172 17264
rect 5224 17252 5230 17264
rect 5353 17255 5411 17261
rect 5353 17252 5365 17255
rect 5224 17224 5365 17252
rect 5224 17212 5230 17224
rect 5353 17221 5365 17224
rect 5399 17221 5411 17255
rect 8386 17252 8392 17264
rect 5353 17215 5411 17221
rect 6656 17224 8392 17252
rect 6656 17184 6684 17224
rect 8386 17212 8392 17224
rect 8444 17252 8450 17264
rect 9122 17252 9128 17264
rect 8444 17224 9128 17252
rect 8444 17212 8450 17224
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 10502 17252 10508 17264
rect 9324 17224 10508 17252
rect 5092 17156 6684 17184
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 7834 17184 7840 17196
rect 6788 17156 6833 17184
rect 7795 17156 7840 17184
rect 6788 17144 6794 17156
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 9324 17193 9352 17224
rect 10502 17212 10508 17224
rect 10560 17212 10566 17264
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17153 9367 17187
rect 9309 17147 9367 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 9539 17156 10149 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10612 17184 10640 17292
rect 12618 17280 12624 17332
rect 12676 17280 12682 17332
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 15010 17320 15016 17332
rect 12768 17292 15016 17320
rect 12768 17280 12774 17292
rect 15010 17280 15016 17292
rect 15068 17320 15074 17332
rect 16114 17320 16120 17332
rect 15068 17292 16120 17320
rect 15068 17280 15074 17292
rect 16114 17280 16120 17292
rect 16172 17280 16178 17332
rect 18414 17280 18420 17332
rect 18472 17320 18478 17332
rect 19889 17323 19947 17329
rect 19889 17320 19901 17323
rect 18472 17292 19901 17320
rect 18472 17280 18478 17292
rect 19889 17289 19901 17292
rect 19935 17289 19947 17323
rect 19889 17283 19947 17289
rect 10781 17255 10839 17261
rect 10781 17221 10793 17255
rect 10827 17252 10839 17255
rect 11146 17252 11152 17264
rect 10827 17224 11152 17252
rect 10827 17221 10839 17224
rect 10781 17215 10839 17221
rect 11146 17212 11152 17224
rect 11204 17212 11210 17264
rect 12636 17252 12664 17280
rect 12636 17224 12747 17252
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 10612 17156 10977 17184
rect 10137 17147 10195 17153
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 12434 17184 12440 17196
rect 12395 17156 12440 17184
rect 10965 17147 11023 17153
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 12719 17193 12747 17224
rect 12693 17187 12751 17193
rect 12693 17153 12705 17187
rect 12739 17153 12751 17187
rect 14458 17184 14464 17196
rect 14419 17156 14464 17184
rect 12693 17147 12751 17153
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 14645 17187 14703 17193
rect 14645 17153 14657 17187
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 1912 17088 3433 17116
rect 1912 17076 1918 17088
rect 3421 17085 3433 17088
rect 3467 17085 3479 17119
rect 6822 17116 6828 17128
rect 6783 17088 6828 17116
rect 3421 17079 3479 17085
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17116 7711 17119
rect 9125 17119 9183 17125
rect 9125 17116 9137 17119
rect 7699 17088 9137 17116
rect 7699 17085 7711 17088
rect 7653 17079 7711 17085
rect 9125 17085 9137 17088
rect 9171 17116 9183 17119
rect 11054 17116 11060 17128
rect 9171 17088 11060 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11882 17116 11888 17128
rect 11195 17088 11888 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 11882 17076 11888 17088
rect 11940 17076 11946 17128
rect 14660 17116 14688 17147
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 15068 17156 15117 17184
rect 15068 17144 15074 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15286 17184 15292 17196
rect 15247 17156 15292 17184
rect 15105 17147 15163 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 15509 17187 15567 17193
rect 15509 17153 15521 17187
rect 15555 17184 15567 17187
rect 15654 17184 15660 17196
rect 15555 17156 15660 17184
rect 15555 17153 15567 17156
rect 15509 17147 15567 17153
rect 15197 17119 15255 17125
rect 15197 17116 15209 17119
rect 14660 17088 15209 17116
rect 15197 17085 15209 17088
rect 15243 17085 15255 17119
rect 15396 17116 15424 17147
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 15746 17144 15752 17196
rect 15804 17184 15810 17196
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 15804 17156 16037 17184
rect 15804 17144 15810 17156
rect 16025 17153 16037 17156
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17184 16267 17187
rect 16666 17184 16672 17196
rect 16255 17156 16672 17184
rect 16255 17153 16267 17156
rect 16209 17147 16267 17153
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 17494 17184 17500 17196
rect 17455 17156 17500 17184
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 18765 17187 18823 17193
rect 18765 17184 18777 17187
rect 18380 17156 18777 17184
rect 18380 17144 18386 17156
rect 18765 17153 18777 17156
rect 18811 17153 18823 17187
rect 18765 17147 18823 17153
rect 16850 17116 16856 17128
rect 15396 17088 16856 17116
rect 15197 17079 15255 17085
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 18414 17076 18420 17128
rect 18472 17116 18478 17128
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18472 17088 18521 17116
rect 18472 17076 18478 17088
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 5537 17051 5595 17057
rect 5537 17017 5549 17051
rect 5583 17048 5595 17051
rect 9030 17048 9036 17060
rect 5583 17020 9036 17048
rect 5583 17017 5595 17020
rect 5537 17011 5595 17017
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 15102 17008 15108 17060
rect 15160 17048 15166 17060
rect 17681 17051 17739 17057
rect 17681 17048 17693 17051
rect 15160 17020 17693 17048
rect 15160 17008 15166 17020
rect 17681 17017 17693 17020
rect 17727 17048 17739 17051
rect 18138 17048 18144 17060
rect 17727 17020 18144 17048
rect 17727 17017 17739 17020
rect 17681 17011 17739 17017
rect 18138 17008 18144 17020
rect 18196 17008 18202 17060
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 8021 16983 8079 16989
rect 8021 16980 8033 16983
rect 7432 16952 8033 16980
rect 7432 16940 7438 16952
rect 8021 16949 8033 16952
rect 8067 16949 8079 16983
rect 9950 16980 9956 16992
rect 9911 16952 9956 16980
rect 8021 16943 8079 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 13630 16980 13636 16992
rect 12860 16952 13636 16980
rect 12860 16940 12866 16952
rect 13630 16940 13636 16952
rect 13688 16980 13694 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 13688 16952 13829 16980
rect 13688 16940 13694 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 14461 16983 14519 16989
rect 14461 16949 14473 16983
rect 14507 16980 14519 16983
rect 15930 16980 15936 16992
rect 14507 16952 15936 16980
rect 14507 16949 14519 16952
rect 14461 16943 14519 16949
rect 15930 16940 15936 16952
rect 15988 16940 15994 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 16080 16952 16129 16980
rect 16080 16940 16086 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 18524 16980 18552 17079
rect 19242 16980 19248 16992
rect 18524 16952 19248 16980
rect 16117 16943 16175 16949
rect 19242 16940 19248 16952
rect 19300 16940 19306 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 4062 16776 4068 16788
rect 4023 16748 4068 16776
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 8389 16779 8447 16785
rect 8389 16776 8401 16779
rect 6880 16748 8401 16776
rect 6880 16736 6886 16748
rect 8389 16745 8401 16748
rect 8435 16776 8447 16779
rect 9398 16776 9404 16788
rect 8435 16748 9404 16776
rect 8435 16745 8447 16748
rect 8389 16739 8447 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 11146 16776 11152 16788
rect 11107 16748 11152 16776
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 15013 16779 15071 16785
rect 15013 16745 15025 16779
rect 15059 16776 15071 16779
rect 15286 16776 15292 16788
rect 15059 16748 15292 16776
rect 15059 16745 15071 16748
rect 15013 16739 15071 16745
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15933 16779 15991 16785
rect 15933 16745 15945 16779
rect 15979 16776 15991 16779
rect 16114 16776 16120 16788
rect 15979 16748 16120 16776
rect 15979 16745 15991 16748
rect 15933 16739 15991 16745
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 18322 16776 18328 16788
rect 18283 16748 18328 16776
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 12897 16711 12955 16717
rect 12897 16708 12909 16711
rect 11808 16680 12909 16708
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16609 7067 16643
rect 9122 16640 9128 16652
rect 9083 16612 9128 16640
rect 7009 16603 7067 16609
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16572 4307 16575
rect 5350 16572 5356 16584
rect 4295 16544 5356 16572
rect 4295 16541 4307 16544
rect 4249 16535 4307 16541
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 6549 16575 6607 16581
rect 6549 16572 6561 16575
rect 6052 16544 6561 16572
rect 6052 16532 6058 16544
rect 6549 16541 6561 16544
rect 6595 16541 6607 16575
rect 6549 16535 6607 16541
rect 7024 16572 7052 16603
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 11808 16649 11836 16680
rect 12897 16677 12909 16680
rect 12943 16677 12955 16711
rect 12897 16671 12955 16677
rect 15194 16668 15200 16720
rect 15252 16708 15258 16720
rect 16485 16711 16543 16717
rect 16485 16708 16497 16711
rect 15252 16680 16497 16708
rect 15252 16668 15258 16680
rect 16485 16677 16497 16680
rect 16531 16677 16543 16711
rect 18506 16708 18512 16720
rect 16485 16671 16543 16677
rect 17604 16680 18512 16708
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 12158 16640 12164 16652
rect 11940 16612 12164 16640
rect 11940 16600 11946 16612
rect 12158 16600 12164 16612
rect 12216 16640 12222 16652
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 12216 16612 12449 16640
rect 12216 16600 12222 16612
rect 12437 16609 12449 16612
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15562 16640 15568 16652
rect 14967 16612 15424 16640
rect 15523 16612 15568 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 8202 16572 8208 16584
rect 7024 16544 8208 16572
rect 6365 16439 6423 16445
rect 6365 16405 6377 16439
rect 6411 16436 6423 16439
rect 7024 16436 7052 16544
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 9392 16575 9450 16581
rect 9392 16541 9404 16575
rect 9438 16572 9450 16575
rect 9950 16572 9956 16584
rect 9438 16544 9956 16572
rect 9438 16541 9450 16544
rect 9392 16535 9450 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 10980 16544 12541 16572
rect 7282 16513 7288 16516
rect 7276 16467 7288 16513
rect 7340 16504 7346 16516
rect 7340 16476 7376 16504
rect 7282 16464 7288 16467
rect 7340 16464 7346 16476
rect 10980 16448 11008 16544
rect 12529 16541 12541 16544
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 12710 16532 12716 16584
rect 12768 16572 12774 16584
rect 13357 16575 13415 16581
rect 13357 16572 13369 16575
rect 12768 16544 13369 16572
rect 12768 16532 12774 16544
rect 13357 16541 13369 16544
rect 13403 16541 13415 16575
rect 13357 16535 13415 16541
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 14829 16575 14887 16581
rect 13504 16544 13549 16572
rect 13504 16532 13510 16544
rect 14829 16541 14841 16575
rect 14875 16541 14887 16575
rect 15396 16572 15424 16612
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 17604 16649 17632 16680
rect 18506 16668 18512 16680
rect 18564 16708 18570 16720
rect 19058 16708 19064 16720
rect 18564 16680 19064 16708
rect 18564 16668 18570 16680
rect 19058 16668 19064 16680
rect 19116 16668 19122 16720
rect 17589 16643 17647 16649
rect 16684 16612 17540 16640
rect 15396 16544 15700 16572
rect 14829 16535 14887 16541
rect 11517 16507 11575 16513
rect 11517 16473 11529 16507
rect 11563 16504 11575 16507
rect 11790 16504 11796 16516
rect 11563 16476 11796 16504
rect 11563 16473 11575 16476
rect 11517 16467 11575 16473
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 13538 16464 13544 16516
rect 13596 16504 13602 16516
rect 14844 16504 14872 16535
rect 13596 16476 14872 16504
rect 15105 16507 15163 16513
rect 13596 16464 13602 16476
rect 15105 16473 15117 16507
rect 15151 16504 15163 16507
rect 15470 16504 15476 16516
rect 15151 16476 15476 16504
rect 15151 16473 15163 16476
rect 15105 16467 15163 16473
rect 15470 16464 15476 16476
rect 15528 16464 15534 16516
rect 15672 16504 15700 16544
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 16390 16572 16396 16584
rect 15804 16544 15849 16572
rect 16351 16544 16396 16572
rect 15804 16532 15810 16544
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 16482 16532 16488 16584
rect 16540 16572 16546 16584
rect 16577 16575 16635 16581
rect 16577 16572 16589 16575
rect 16540 16544 16589 16572
rect 16540 16532 16546 16544
rect 16577 16541 16589 16544
rect 16623 16541 16635 16575
rect 16577 16535 16635 16541
rect 16408 16504 16436 16532
rect 16684 16504 16712 16612
rect 17218 16532 17224 16584
rect 17276 16532 17282 16584
rect 17512 16572 17540 16612
rect 17589 16609 17601 16643
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16609 17739 16643
rect 17681 16603 17739 16609
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16640 17923 16643
rect 18046 16640 18052 16652
rect 17911 16612 18052 16640
rect 17911 16609 17923 16612
rect 17865 16603 17923 16609
rect 17696 16572 17724 16603
rect 18046 16600 18052 16612
rect 18104 16600 18110 16652
rect 17512 16544 17724 16572
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16572 18567 16575
rect 18782 16572 18788 16584
rect 18555 16544 18788 16572
rect 18555 16541 18567 16544
rect 18509 16535 18567 16541
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 15672 16476 16436 16504
rect 16500 16476 16712 16504
rect 17236 16504 17264 16532
rect 17586 16504 17592 16516
rect 17236 16476 17592 16504
rect 6411 16408 7052 16436
rect 10505 16439 10563 16445
rect 6411 16405 6423 16408
rect 6365 16399 6423 16405
rect 10505 16405 10517 16439
rect 10551 16436 10563 16439
rect 10962 16436 10968 16448
rect 10551 16408 10968 16436
rect 10551 16405 10563 16408
rect 10505 16399 10563 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 11609 16439 11667 16445
rect 11609 16405 11621 16439
rect 11655 16436 11667 16439
rect 12250 16436 12256 16448
rect 11655 16408 12256 16436
rect 11655 16405 11667 16408
rect 11609 16399 11667 16405
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 16500 16436 16528 16476
rect 17586 16464 17592 16476
rect 17644 16464 17650 16516
rect 15712 16408 16528 16436
rect 17221 16439 17279 16445
rect 15712 16396 15718 16408
rect 17221 16405 17233 16439
rect 17267 16436 17279 16439
rect 17310 16436 17316 16448
rect 17267 16408 17316 16436
rect 17267 16405 17279 16408
rect 17221 16399 17279 16405
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16232 7251 16235
rect 7282 16232 7288 16244
rect 7239 16204 7288 16232
rect 7239 16201 7251 16204
rect 7193 16195 7251 16201
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 10778 16232 10784 16244
rect 10367 16204 10784 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 10778 16192 10784 16204
rect 10836 16232 10842 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10836 16204 11069 16232
rect 10836 16192 10842 16204
rect 11057 16201 11069 16204
rect 11103 16232 11115 16235
rect 11514 16232 11520 16244
rect 11103 16204 11520 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 14921 16235 14979 16241
rect 14921 16201 14933 16235
rect 14967 16232 14979 16235
rect 15378 16232 15384 16244
rect 14967 16204 15384 16232
rect 14967 16201 14979 16204
rect 14921 16195 14979 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 15562 16192 15568 16244
rect 15620 16232 15626 16244
rect 16298 16232 16304 16244
rect 15620 16204 16304 16232
rect 15620 16192 15626 16204
rect 16298 16192 16304 16204
rect 16356 16232 16362 16244
rect 17221 16235 17279 16241
rect 16356 16204 17172 16232
rect 16356 16192 16362 16204
rect 10962 16164 10968 16176
rect 10923 16136 10968 16164
rect 10962 16124 10968 16136
rect 11020 16164 11026 16176
rect 12618 16164 12624 16176
rect 11020 16136 12624 16164
rect 11020 16124 11026 16136
rect 12618 16124 12624 16136
rect 12676 16164 12682 16176
rect 12676 16136 12848 16164
rect 12676 16124 12682 16136
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 9033 16099 9091 16105
rect 9033 16096 9045 16099
rect 8812 16068 9045 16096
rect 8812 16056 8818 16068
rect 9033 16065 9045 16068
rect 9079 16065 9091 16099
rect 9033 16059 9091 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16096 10195 16099
rect 10318 16096 10324 16108
rect 10183 16068 10324 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 10870 16096 10876 16108
rect 10459 16068 10876 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 10870 16056 10876 16068
rect 10928 16096 10934 16108
rect 11698 16096 11704 16108
rect 10928 16068 11704 16096
rect 10928 16056 10934 16068
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 11882 16096 11888 16108
rect 11843 16068 11888 16096
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16065 12035 16099
rect 12250 16096 12256 16108
rect 12211 16068 12256 16096
rect 11977 16059 12035 16065
rect 11992 16028 12020 16059
rect 12250 16056 12256 16068
rect 12308 16056 12314 16108
rect 12710 16096 12716 16108
rect 12671 16068 12716 16096
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 12820 16105 12848 16136
rect 15470 16124 15476 16176
rect 15528 16164 15534 16176
rect 15933 16167 15991 16173
rect 15933 16164 15945 16167
rect 15528 16136 15945 16164
rect 15528 16124 15534 16136
rect 15933 16133 15945 16136
rect 15979 16164 15991 16167
rect 16482 16164 16488 16176
rect 15979 16136 16488 16164
rect 15979 16133 15991 16136
rect 15933 16127 15991 16133
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 16853 16167 16911 16173
rect 16853 16133 16865 16167
rect 16899 16133 16911 16167
rect 16853 16127 16911 16133
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 12894 16056 12900 16108
rect 12952 16096 12958 16108
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 12952 16068 13737 16096
rect 12952 16056 12958 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 15102 16096 15108 16108
rect 15063 16068 15108 16096
rect 13725 16059 13783 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 15286 16096 15292 16108
rect 15247 16068 15292 16096
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15838 16096 15844 16108
rect 15799 16068 15844 16096
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 16868 16096 16896 16127
rect 17034 16124 17040 16176
rect 17092 16173 17098 16176
rect 17092 16167 17111 16173
rect 17099 16133 17111 16167
rect 17144 16164 17172 16204
rect 17221 16201 17233 16235
rect 17267 16232 17279 16235
rect 17586 16232 17592 16244
rect 17267 16204 17592 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 19058 16232 19064 16244
rect 19019 16204 19064 16232
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 17144 16136 17356 16164
rect 17092 16127 17111 16133
rect 17092 16124 17098 16127
rect 17218 16096 17224 16108
rect 16868 16068 17224 16096
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 17328 16096 17356 16136
rect 17402 16124 17408 16176
rect 17460 16164 17466 16176
rect 18414 16164 18420 16176
rect 17460 16136 18420 16164
rect 17460 16124 17466 16136
rect 18414 16124 18420 16136
rect 18472 16124 18478 16176
rect 18506 16124 18512 16176
rect 18564 16164 18570 16176
rect 22278 16164 22284 16176
rect 18564 16136 22284 16164
rect 18564 16124 18570 16136
rect 22278 16124 22284 16136
rect 22336 16124 22342 16176
rect 17328 16068 17540 16096
rect 12728 16028 12756 16056
rect 13538 16028 13544 16040
rect 10152 16000 12020 16028
rect 12084 16000 12756 16028
rect 13499 16000 13544 16028
rect 10152 15969 10180 16000
rect 10137 15963 10195 15969
rect 10137 15929 10149 15963
rect 10183 15929 10195 15963
rect 10137 15923 10195 15929
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 11330 15960 11336 15972
rect 10376 15932 11336 15960
rect 10376 15920 10382 15932
rect 11330 15920 11336 15932
rect 11388 15960 11394 15972
rect 12084 15960 12112 16000
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 15378 16028 15384 16040
rect 15339 16000 15384 16028
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 16206 16028 16212 16040
rect 16167 16000 16212 16028
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 17512 16028 17540 16068
rect 18782 16056 18788 16108
rect 18840 16096 18846 16108
rect 18969 16099 19027 16105
rect 18969 16096 18981 16099
rect 18840 16068 18981 16096
rect 18840 16056 18846 16068
rect 18969 16065 18981 16068
rect 19015 16065 19027 16099
rect 18969 16059 19027 16065
rect 17681 16031 17739 16037
rect 17681 16028 17693 16031
rect 17512 16000 17693 16028
rect 17681 15997 17693 16000
rect 17727 15997 17739 16031
rect 17681 15991 17739 15997
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 16028 18015 16031
rect 19610 16028 19616 16040
rect 18003 16000 19616 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 11388 15932 12112 15960
rect 11388 15920 11394 15932
rect 9217 15895 9275 15901
rect 9217 15861 9229 15895
rect 9263 15892 9275 15895
rect 9306 15892 9312 15904
rect 9263 15864 9312 15892
rect 9263 15861 9275 15864
rect 9217 15855 9275 15861
rect 9306 15852 9312 15864
rect 9364 15892 9370 15904
rect 11422 15892 11428 15904
rect 9364 15864 11428 15892
rect 9364 15852 9370 15864
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 11698 15892 11704 15904
rect 11659 15864 11704 15892
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 12802 15892 12808 15904
rect 12763 15864 12808 15892
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 13081 15895 13139 15901
rect 13081 15892 13093 15895
rect 13044 15864 13093 15892
rect 13044 15852 13050 15864
rect 13081 15861 13093 15864
rect 13127 15861 13139 15895
rect 13906 15892 13912 15904
rect 13867 15864 13912 15892
rect 13081 15855 13139 15861
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 16022 15892 16028 15904
rect 14608 15864 16028 15892
rect 14608 15852 14614 15864
rect 16022 15852 16028 15864
rect 16080 15892 16086 15904
rect 16117 15895 16175 15901
rect 16117 15892 16129 15895
rect 16080 15864 16129 15892
rect 16080 15852 16086 15864
rect 16117 15861 16129 15864
rect 16163 15861 16175 15895
rect 16298 15892 16304 15904
rect 16259 15864 16304 15892
rect 16117 15855 16175 15861
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 16942 15892 16948 15904
rect 16448 15864 16948 15892
rect 16448 15852 16454 15864
rect 16942 15852 16948 15864
rect 17000 15892 17006 15904
rect 17037 15895 17095 15901
rect 17037 15892 17049 15895
rect 17000 15864 17049 15892
rect 17000 15852 17006 15864
rect 17037 15861 17049 15864
rect 17083 15892 17095 15895
rect 18064 15892 18092 16000
rect 19610 15988 19616 16000
rect 19668 15988 19674 16040
rect 17083 15864 18092 15892
rect 17083 15861 17095 15864
rect 17037 15855 17095 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 11333 15691 11391 15697
rect 11333 15657 11345 15691
rect 11379 15688 11391 15691
rect 11882 15688 11888 15700
rect 11379 15660 11888 15688
rect 11379 15657 11391 15660
rect 11333 15651 11391 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 14829 15691 14887 15697
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 16206 15688 16212 15700
rect 14875 15660 16212 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17218 15648 17224 15700
rect 17276 15688 17282 15700
rect 17678 15688 17684 15700
rect 17276 15660 17684 15688
rect 17276 15648 17282 15660
rect 17678 15648 17684 15660
rect 17736 15688 17742 15700
rect 18782 15688 18788 15700
rect 17736 15660 18788 15688
rect 17736 15648 17742 15660
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 10778 15580 10784 15632
rect 10836 15620 10842 15632
rect 12618 15620 12624 15632
rect 10836 15592 11744 15620
rect 12579 15592 12624 15620
rect 10836 15580 10842 15592
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 8938 15552 8944 15564
rect 8812 15524 8944 15552
rect 8812 15512 8818 15524
rect 8938 15512 8944 15524
rect 8996 15552 9002 15564
rect 9309 15555 9367 15561
rect 9309 15552 9321 15555
rect 8996 15524 9321 15552
rect 8996 15512 9002 15524
rect 9309 15521 9321 15524
rect 9355 15552 9367 15555
rect 11238 15552 11244 15564
rect 9355 15524 11244 15552
rect 9355 15521 9367 15524
rect 9309 15515 9367 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 11716 15561 11744 15592
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 15378 15620 15384 15632
rect 15291 15592 15384 15620
rect 15378 15580 15384 15592
rect 15436 15620 15442 15632
rect 16574 15620 16580 15632
rect 15436 15592 16580 15620
rect 15436 15580 15442 15592
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 11517 15555 11575 15561
rect 11517 15552 11529 15555
rect 11388 15524 11529 15552
rect 11388 15512 11394 15524
rect 11517 15521 11529 15524
rect 11563 15521 11575 15555
rect 11517 15515 11575 15521
rect 11692 15555 11750 15561
rect 11692 15521 11704 15555
rect 11738 15521 11750 15555
rect 11692 15515 11750 15521
rect 11790 15512 11796 15564
rect 11848 15552 11854 15564
rect 11848 15524 11893 15552
rect 11848 15512 11854 15524
rect 13538 15512 13544 15564
rect 13596 15552 13602 15564
rect 15473 15555 15531 15561
rect 15473 15552 15485 15555
rect 13596 15524 15485 15552
rect 13596 15512 13602 15524
rect 15473 15521 15485 15524
rect 15519 15521 15531 15555
rect 15473 15515 15531 15521
rect 16298 15512 16304 15564
rect 16356 15552 16362 15564
rect 16853 15555 16911 15561
rect 16853 15552 16865 15555
rect 16356 15524 16865 15552
rect 16356 15512 16362 15524
rect 16853 15521 16865 15524
rect 16899 15552 16911 15555
rect 16899 15524 17540 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 9088 15456 9137 15484
rect 9088 15444 9094 15456
rect 9125 15453 9137 15456
rect 9171 15484 9183 15487
rect 9214 15484 9220 15496
rect 9171 15456 9220 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 10008 15456 10057 15484
rect 10008 15444 10014 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 10045 15447 10103 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 11598 15487 11656 15493
rect 11598 15453 11610 15487
rect 11644 15453 11656 15487
rect 11598 15447 11656 15453
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11624 15348 11652 15447
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 12032 15456 12909 15484
rect 12032 15444 12038 15456
rect 12897 15453 12909 15456
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13078 15484 13084 15496
rect 13035 15456 13084 15484
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 15010 15487 15068 15493
rect 15010 15453 15022 15487
rect 15056 15484 15068 15487
rect 15378 15484 15384 15496
rect 15056 15456 15384 15484
rect 15056 15453 15068 15456
rect 15010 15447 15068 15453
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15654 15444 15660 15496
rect 15712 15484 15718 15496
rect 16485 15487 16543 15493
rect 16485 15484 16497 15487
rect 15712 15456 16497 15484
rect 15712 15444 15718 15456
rect 16485 15453 16497 15456
rect 16531 15453 16543 15487
rect 16485 15447 16543 15453
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 16758 15484 16764 15496
rect 16623 15456 16764 15484
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 16758 15444 16764 15456
rect 16816 15444 16822 15496
rect 16942 15484 16948 15496
rect 16903 15456 16948 15484
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17402 15484 17408 15496
rect 17363 15456 17408 15484
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 17512 15484 17540 15524
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 17512 15456 19441 15484
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19610 15484 19616 15496
rect 19571 15456 19616 15484
rect 19429 15447 19487 15453
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 12802 15416 12808 15428
rect 12763 15388 12808 15416
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 16209 15419 16267 15425
rect 16209 15385 16221 15419
rect 16255 15416 16267 15419
rect 17218 15416 17224 15428
rect 16255 15388 17224 15416
rect 16255 15385 16267 15388
rect 16209 15379 16267 15385
rect 17218 15376 17224 15388
rect 17276 15376 17282 15428
rect 17672 15419 17730 15425
rect 17672 15385 17684 15419
rect 17718 15416 17730 15419
rect 17954 15416 17960 15428
rect 17718 15388 17960 15416
rect 17718 15385 17730 15388
rect 17672 15379 17730 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 19521 15419 19579 15425
rect 19521 15416 19533 15419
rect 18064 15388 19533 15416
rect 10928 15320 11652 15348
rect 13173 15351 13231 15357
rect 10928 15308 10934 15320
rect 13173 15317 13185 15351
rect 13219 15348 13231 15351
rect 13262 15348 13268 15360
rect 13219 15320 13268 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 15013 15351 15071 15357
rect 15013 15317 15025 15351
rect 15059 15348 15071 15351
rect 15194 15348 15200 15360
rect 15059 15320 15200 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 16669 15351 16727 15357
rect 16669 15317 16681 15351
rect 16715 15348 16727 15351
rect 18064 15348 18092 15388
rect 19521 15385 19533 15388
rect 19567 15385 19579 15419
rect 19521 15379 19579 15385
rect 16715 15320 18092 15348
rect 16715 15317 16727 15320
rect 16669 15311 16727 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 9950 15144 9956 15156
rect 9815 15116 9956 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 10410 15144 10416 15156
rect 10371 15116 10416 15144
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 11701 15147 11759 15153
rect 11701 15113 11713 15147
rect 11747 15144 11759 15147
rect 11882 15144 11888 15156
rect 11747 15116 11888 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 13357 15147 13415 15153
rect 12308 15116 13308 15144
rect 12308 15104 12314 15116
rect 8386 15008 8392 15020
rect 8347 14980 8392 15008
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 8656 15011 8714 15017
rect 8656 14977 8668 15011
rect 8702 15008 8714 15011
rect 9122 15008 9128 15020
rect 8702 14980 9128 15008
rect 8702 14977 8714 14980
rect 8656 14971 8714 14977
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 10318 14968 10324 15020
rect 10376 15017 10382 15020
rect 10376 15011 10412 15017
rect 10400 14977 10412 15011
rect 10376 14971 10412 14977
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 15008 10931 15011
rect 11698 15008 11704 15020
rect 10919 14980 11704 15008
rect 10919 14977 10931 14980
rect 10873 14971 10931 14977
rect 10376 14968 10382 14971
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 11848 14980 12081 15008
rect 11848 14968 11854 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 15008 12219 15011
rect 12526 15008 12532 15020
rect 12207 14980 12532 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 12526 14968 12532 14980
rect 12584 15008 12590 15020
rect 12986 15008 12992 15020
rect 12584 14980 12992 15008
rect 12584 14968 12590 14980
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 13078 14968 13084 15020
rect 13136 15008 13142 15020
rect 13136 14980 13181 15008
rect 13136 14968 13142 14980
rect 13280 14940 13308 15116
rect 13357 15113 13369 15147
rect 13403 15113 13415 15147
rect 13357 15107 13415 15113
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15102 15144 15108 15156
rect 15059 15116 15108 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 13372 15008 13400 15107
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 15804 15116 17233 15144
rect 15804 15104 15810 15116
rect 17221 15113 17233 15116
rect 17267 15113 17279 15147
rect 17221 15107 17279 15113
rect 16574 15036 16580 15088
rect 16632 15076 16638 15088
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 16632 15048 17049 15076
rect 16632 15036 16638 15048
rect 17037 15045 17049 15048
rect 17083 15045 17095 15079
rect 17037 15039 17095 15045
rect 13538 15008 13544 15020
rect 13372 14980 13544 15008
rect 13538 14968 13544 14980
rect 13596 15008 13602 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13596 14980 14197 15008
rect 13596 14968 13602 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14274 14968 14280 15020
rect 14332 15008 14338 15020
rect 14458 15008 14464 15020
rect 14332 14980 14377 15008
rect 14419 14980 14464 15008
rect 14332 14968 14338 14980
rect 14458 14968 14464 14980
rect 14516 14968 14522 15020
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 15289 15011 15347 15017
rect 14608 14980 14653 15008
rect 14608 14968 14614 14980
rect 15289 14977 15301 15011
rect 15335 15008 15347 15011
rect 16390 15008 16396 15020
rect 15335 14980 16396 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 16482 14968 16488 15020
rect 16540 15008 16546 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16540 14980 16865 15008
rect 16540 14968 16546 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 17678 15008 17684 15020
rect 17639 14980 17684 15008
rect 16853 14971 16911 14977
rect 17678 14968 17684 14980
rect 17736 14968 17742 15020
rect 13722 14940 13728 14952
rect 13280 14912 13728 14940
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 10042 14832 10048 14884
rect 10100 14872 10106 14884
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 10100 14844 10793 14872
rect 10100 14832 10106 14844
rect 10781 14841 10793 14844
rect 10827 14872 10839 14875
rect 12618 14872 12624 14884
rect 10827 14844 12624 14872
rect 10827 14841 10839 14844
rect 10781 14835 10839 14841
rect 12618 14832 12624 14844
rect 12676 14832 12682 14884
rect 14292 14872 14320 14968
rect 15194 14940 15200 14952
rect 15155 14912 15200 14940
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 15378 14940 15384 14952
rect 15339 14912 15384 14940
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 15473 14943 15531 14949
rect 15473 14909 15485 14943
rect 15519 14940 15531 14943
rect 15838 14940 15844 14952
rect 15519 14912 15844 14940
rect 15519 14909 15531 14912
rect 15473 14903 15531 14909
rect 15286 14872 15292 14884
rect 14292 14844 15292 14872
rect 15286 14832 15292 14844
rect 15344 14872 15350 14884
rect 15488 14872 15516 14903
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 17770 14900 17776 14952
rect 17828 14940 17834 14952
rect 17957 14943 18015 14949
rect 17957 14940 17969 14943
rect 17828 14912 17969 14940
rect 17828 14900 17834 14912
rect 17957 14909 17969 14912
rect 18003 14909 18015 14943
rect 17957 14903 18015 14909
rect 15344 14844 15516 14872
rect 15344 14832 15350 14844
rect 16758 14832 16764 14884
rect 16816 14872 16822 14884
rect 18230 14872 18236 14884
rect 16816 14844 18236 14872
rect 16816 14832 16822 14844
rect 18230 14832 18236 14844
rect 18288 14832 18294 14884
rect 10226 14804 10232 14816
rect 10187 14776 10232 14804
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 12342 14804 12348 14816
rect 12303 14776 12348 14804
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 13170 14804 13176 14816
rect 13131 14776 13176 14804
rect 13170 14764 13176 14776
rect 13228 14804 13234 14816
rect 13814 14804 13820 14816
rect 13228 14776 13820 14804
rect 13228 14764 13234 14776
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 13998 14804 14004 14816
rect 13959 14776 14004 14804
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 17770 14804 17776 14816
rect 15436 14776 17776 14804
rect 15436 14764 15442 14776
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 9122 14600 9128 14612
rect 9083 14572 9128 14600
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 10870 14600 10876 14612
rect 10831 14572 10876 14600
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 11885 14603 11943 14609
rect 11885 14569 11897 14603
rect 11931 14600 11943 14603
rect 12158 14600 12164 14612
rect 11931 14572 12164 14600
rect 11931 14569 11943 14572
rect 11885 14563 11943 14569
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 12894 14600 12900 14612
rect 12667 14572 12900 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 13906 14600 13912 14612
rect 13679 14572 13912 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14458 14600 14464 14612
rect 14419 14572 14464 14600
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 15562 14560 15568 14612
rect 15620 14600 15626 14612
rect 17037 14603 17095 14609
rect 17037 14600 17049 14603
rect 15620 14572 17049 14600
rect 15620 14560 15626 14572
rect 17037 14569 17049 14572
rect 17083 14569 17095 14603
rect 17037 14563 17095 14569
rect 17129 14603 17187 14609
rect 17129 14569 17141 14603
rect 17175 14600 17187 14603
rect 17678 14600 17684 14612
rect 17175 14572 17684 14600
rect 17175 14569 17187 14572
rect 17129 14563 17187 14569
rect 17678 14560 17684 14572
rect 17736 14560 17742 14612
rect 17954 14600 17960 14612
rect 17915 14572 17960 14600
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 9306 14532 9312 14544
rect 2746 14504 9312 14532
rect 1946 14424 1952 14476
rect 2004 14464 2010 14476
rect 2746 14464 2774 14504
rect 9306 14492 9312 14504
rect 9364 14492 9370 14544
rect 10226 14464 10232 14476
rect 2004 14436 2774 14464
rect 9140 14436 10232 14464
rect 2004 14424 2010 14436
rect 9140 14405 9168 14436
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 10376 14436 11069 14464
rect 10376 14424 10382 14436
rect 11057 14433 11069 14436
rect 11103 14433 11115 14467
rect 12544 14464 12572 14560
rect 13998 14492 14004 14544
rect 14056 14532 14062 14544
rect 17310 14532 17316 14544
rect 14056 14504 17316 14532
rect 14056 14492 14062 14504
rect 17310 14492 17316 14504
rect 17368 14532 17374 14544
rect 17865 14535 17923 14541
rect 17865 14532 17877 14535
rect 17368 14504 17877 14532
rect 17368 14492 17374 14504
rect 17865 14501 17877 14504
rect 17911 14501 17923 14535
rect 17865 14495 17923 14501
rect 11057 14427 11115 14433
rect 11716 14436 12572 14464
rect 12713 14467 12771 14473
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14365 9183 14399
rect 9306 14396 9312 14408
rect 9267 14368 9312 14396
rect 9125 14359 9183 14365
rect 9306 14356 9312 14368
rect 9364 14396 9370 14408
rect 10502 14396 10508 14408
rect 9364 14368 10508 14396
rect 9364 14356 9370 14368
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 10778 14396 10784 14408
rect 10739 14368 10784 14396
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11716 14405 11744 14436
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 12802 14464 12808 14476
rect 12759 14436 12808 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 12802 14424 12808 14436
rect 12860 14464 12866 14476
rect 13170 14464 13176 14476
rect 12860 14436 13176 14464
rect 12860 14424 12866 14436
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 18046 14464 18052 14476
rect 13596 14436 17356 14464
rect 18007 14436 18052 14464
rect 13596 14424 13602 14436
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 11057 14331 11115 14337
rect 11057 14297 11069 14331
rect 11103 14328 11115 14331
rect 11532 14328 11560 14359
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12437 14399 12495 14405
rect 12437 14396 12449 14399
rect 11848 14368 12449 14396
rect 11848 14356 11854 14368
rect 12437 14365 12449 14368
rect 12483 14396 12495 14399
rect 13078 14396 13084 14408
rect 12483 14368 13084 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 11103 14300 11560 14328
rect 13372 14328 13400 14359
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 13722 14396 13728 14408
rect 13504 14368 13549 14396
rect 13683 14368 13728 14396
rect 13504 14356 13510 14368
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 14366 14396 14372 14408
rect 14327 14368 14372 14396
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 15010 14396 15016 14408
rect 14971 14368 15016 14396
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 14384 14328 14412 14356
rect 13372 14300 14412 14328
rect 16868 14328 16896 14359
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17328 14405 17356 14436
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 18141 14467 18199 14473
rect 18141 14433 18153 14467
rect 18187 14464 18199 14467
rect 18230 14464 18236 14476
rect 18187 14436 18236 14464
rect 18187 14433 18199 14436
rect 18141 14427 18199 14433
rect 18230 14424 18236 14436
rect 18288 14424 18294 14476
rect 17313 14399 17371 14405
rect 17000 14368 17045 14396
rect 17000 14356 17006 14368
rect 17313 14365 17325 14399
rect 17359 14365 17371 14399
rect 17770 14396 17776 14408
rect 17731 14368 17776 14396
rect 17313 14359 17371 14365
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14396 19671 14399
rect 20070 14396 20076 14408
rect 19659 14368 20076 14396
rect 19659 14365 19671 14368
rect 19613 14359 19671 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 18598 14328 18604 14340
rect 16868 14300 18604 14328
rect 11103 14297 11115 14300
rect 11057 14291 11115 14297
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 13170 14260 13176 14272
rect 13131 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 16577 14263 16635 14269
rect 16577 14260 16589 14263
rect 16540 14232 16589 14260
rect 16540 14220 16546 14232
rect 16577 14229 16589 14232
rect 16623 14229 16635 14263
rect 19426 14260 19432 14272
rect 19387 14232 19432 14260
rect 16577 14223 16635 14229
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9858 14016 9864 14068
rect 9916 14056 9922 14068
rect 10410 14056 10416 14068
rect 9916 14028 10416 14056
rect 9916 14016 9922 14028
rect 10410 14016 10416 14028
rect 10468 14056 10474 14068
rect 12253 14059 12311 14065
rect 12253 14056 12265 14059
rect 10468 14028 12265 14056
rect 10468 14016 10474 14028
rect 12253 14025 12265 14028
rect 12299 14025 12311 14059
rect 12253 14019 12311 14025
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 15068 14028 15117 14056
rect 15068 14016 15074 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 15473 14059 15531 14065
rect 15473 14025 15485 14059
rect 15519 14056 15531 14059
rect 15562 14056 15568 14068
rect 15519 14028 15568 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 15562 14016 15568 14028
rect 15620 14056 15626 14068
rect 18509 14059 18567 14065
rect 18509 14056 18521 14059
rect 15620 14028 18521 14056
rect 15620 14016 15626 14028
rect 18509 14025 18521 14028
rect 18555 14025 18567 14059
rect 18509 14019 18567 14025
rect 9585 13991 9643 13997
rect 9585 13957 9597 13991
rect 9631 13988 9643 13991
rect 10870 13988 10876 14000
rect 9631 13960 10876 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 12802 13988 12808 14000
rect 12636 13960 12808 13988
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 1946 13920 1952 13932
rect 1627 13892 1952 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 9784 13852 9812 13883
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10505 13923 10563 13929
rect 9916 13892 9961 13920
rect 9916 13880 9922 13892
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 10962 13920 10968 13932
rect 10551 13892 10968 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10520 13852 10548 13883
rect 10962 13880 10968 13892
rect 11020 13920 11026 13932
rect 11790 13920 11796 13932
rect 11020 13892 11796 13920
rect 11020 13880 11026 13892
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 12250 13923 12308 13929
rect 12250 13889 12262 13923
rect 12296 13920 12308 13923
rect 12636 13920 12664 13960
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 16301 13991 16359 13997
rect 16301 13988 16313 13991
rect 15580 13960 16313 13988
rect 15580 13932 15608 13960
rect 16301 13957 16313 13960
rect 16347 13988 16359 13991
rect 17034 13988 17040 14000
rect 16347 13960 17040 13988
rect 16347 13957 16359 13960
rect 16301 13951 16359 13957
rect 17034 13948 17040 13960
rect 17092 13948 17098 14000
rect 12296 13892 12664 13920
rect 12713 13923 12771 13929
rect 12296 13889 12308 13892
rect 12250 13883 12308 13889
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 13170 13920 13176 13932
rect 12759 13892 13176 13920
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 13538 13920 13544 13932
rect 13499 13892 13544 13920
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 13814 13920 13820 13932
rect 13775 13892 13820 13920
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 15286 13920 15292 13932
rect 15247 13892 15292 13920
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16942 13920 16948 13932
rect 16163 13892 16948 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17126 13920 17132 13932
rect 17087 13892 17132 13920
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 17218 13880 17224 13932
rect 17276 13920 17282 13932
rect 17385 13923 17443 13929
rect 17385 13920 17397 13923
rect 17276 13892 17397 13920
rect 17276 13880 17282 13892
rect 17385 13889 17397 13892
rect 17431 13889 17443 13923
rect 17385 13883 17443 13889
rect 9784 13824 10548 13852
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 12342 13852 12348 13864
rect 10643 13824 12348 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12618 13784 12624 13796
rect 12579 13756 12624 13784
rect 12618 13744 12624 13756
rect 12676 13744 12682 13796
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 9858 13716 9864 13728
rect 9631 13688 9864 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10836 13688 10885 13716
rect 10836 13676 10842 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 10873 13679 10931 13685
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 12069 13719 12127 13725
rect 12069 13716 12081 13719
rect 11664 13688 12081 13716
rect 11664 13676 11670 13688
rect 12069 13685 12081 13688
rect 12115 13685 12127 13719
rect 12069 13679 12127 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 10962 13512 10968 13524
rect 10919 13484 10968 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 13538 13472 13544 13524
rect 13596 13512 13602 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13596 13484 13645 13512
rect 13596 13472 13602 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 15105 13515 15163 13521
rect 15105 13512 15117 13515
rect 14424 13484 15117 13512
rect 14424 13472 14430 13484
rect 15105 13481 15117 13484
rect 15151 13481 15163 13515
rect 15105 13475 15163 13481
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 17037 13515 17095 13521
rect 17037 13512 17049 13515
rect 17000 13484 17049 13512
rect 17000 13472 17006 13484
rect 17037 13481 17049 13484
rect 17083 13481 17095 13515
rect 17037 13475 17095 13481
rect 8202 13336 8208 13388
rect 8260 13376 8266 13388
rect 9493 13379 9551 13385
rect 9493 13376 9505 13379
rect 8260 13348 9505 13376
rect 8260 13336 8266 13348
rect 9493 13345 9505 13348
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 10560 13348 11836 13376
rect 10560 13336 10566 13348
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11808 13317 11836 13348
rect 14476 13348 15700 13376
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13308 12311 13311
rect 14476 13308 14504 13348
rect 12299 13280 14504 13308
rect 14921 13311 14979 13317
rect 12299 13277 12311 13280
rect 12253 13271 12311 13277
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 15010 13308 15016 13320
rect 14967 13280 15016 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 15672 13317 15700 13348
rect 15930 13317 15936 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 15924 13308 15936 13317
rect 15891 13280 15936 13308
rect 15657 13271 15715 13277
rect 15924 13271 15936 13280
rect 9760 13243 9818 13249
rect 9760 13209 9772 13243
rect 9806 13240 9818 13243
rect 9950 13240 9956 13252
rect 9806 13212 9956 13240
rect 9806 13209 9818 13212
rect 9760 13203 9818 13209
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 11701 13243 11759 13249
rect 11701 13209 11713 13243
rect 11747 13240 11759 13243
rect 12498 13243 12556 13249
rect 12498 13240 12510 13243
rect 11747 13212 12510 13240
rect 11747 13209 11759 13212
rect 11701 13203 11759 13209
rect 12498 13209 12510 13212
rect 12544 13209 12556 13243
rect 14734 13240 14740 13252
rect 14695 13212 14740 13240
rect 12498 13203 12556 13209
rect 14734 13200 14740 13212
rect 14792 13240 14798 13252
rect 15194 13240 15200 13252
rect 14792 13212 15200 13240
rect 14792 13200 14798 13212
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 15672 13240 15700 13271
rect 15930 13268 15936 13271
rect 15988 13268 15994 13320
rect 17126 13240 17132 13252
rect 15672 13212 17132 13240
rect 17126 13200 17132 13212
rect 17184 13200 17190 13252
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 9950 12968 9956 12980
rect 9911 12940 9956 12968
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 10870 12968 10876 12980
rect 10831 12940 10876 12968
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 13265 12971 13323 12977
rect 13265 12937 13277 12971
rect 13311 12968 13323 12971
rect 13446 12968 13452 12980
rect 13311 12940 13452 12968
rect 13311 12937 13323 12940
rect 13265 12931 13323 12937
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 14734 12968 14740 12980
rect 14231 12940 14740 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 15470 12968 15476 12980
rect 15431 12940 15476 12968
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 18598 12968 18604 12980
rect 18559 12940 18604 12968
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 10594 12860 10600 12912
rect 10652 12900 10658 12912
rect 15286 12900 15292 12912
rect 10652 12872 11008 12900
rect 10652 12860 10658 12872
rect 9858 12832 9864 12844
rect 9819 12804 9864 12832
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12832 10103 12835
rect 10502 12832 10508 12844
rect 10091 12804 10508 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 10980 12841 11008 12872
rect 13280 12872 14044 12900
rect 15247 12872 15292 12900
rect 13280 12844 13308 12872
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13262 12832 13268 12844
rect 13219 12804 13268 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 13372 12764 13400 12795
rect 13538 12792 13544 12844
rect 13596 12832 13602 12844
rect 14016 12841 14044 12872
rect 15286 12860 15292 12872
rect 15344 12860 15350 12912
rect 13817 12835 13875 12841
rect 13817 12832 13829 12835
rect 13596 12804 13829 12832
rect 13596 12792 13602 12804
rect 13817 12801 13829 12804
rect 13863 12801 13875 12835
rect 13817 12795 13875 12801
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15010 12832 15016 12844
rect 14875 12804 15016 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 12860 12736 13400 12764
rect 14660 12764 14688 12795
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 15562 12832 15568 12844
rect 15523 12804 15568 12832
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12832 18567 12835
rect 19334 12832 19340 12844
rect 18555 12804 19340 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 19334 12792 19340 12804
rect 19392 12792 19398 12844
rect 38286 12832 38292 12844
rect 38247 12804 38292 12832
rect 38286 12792 38292 12804
rect 38344 12792 38350 12844
rect 16482 12764 16488 12776
rect 14660 12736 16488 12764
rect 12860 12724 12866 12736
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 13722 12656 13728 12708
rect 13780 12696 13786 12708
rect 14737 12699 14795 12705
rect 14737 12696 14749 12699
rect 13780 12668 14749 12696
rect 13780 12656 13786 12668
rect 14737 12665 14749 12668
rect 14783 12665 14795 12699
rect 14737 12659 14795 12665
rect 15289 12699 15347 12705
rect 15289 12665 15301 12699
rect 15335 12696 15347 12699
rect 16574 12696 16580 12708
rect 15335 12668 16580 12696
rect 15335 12665 15347 12668
rect 15289 12659 15347 12665
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 17034 12656 17040 12708
rect 17092 12696 17098 12708
rect 17092 12668 22094 12696
rect 17092 12656 17098 12668
rect 22066 12628 22094 12668
rect 38105 12631 38163 12637
rect 38105 12628 38117 12631
rect 22066 12600 38117 12628
rect 38105 12597 38117 12600
rect 38151 12597 38163 12631
rect 38105 12591 38163 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 17494 12424 17500 12436
rect 17455 12396 17500 12424
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 17313 12359 17371 12365
rect 17313 12356 17325 12359
rect 6604 12328 17325 12356
rect 6604 12316 6610 12328
rect 17313 12325 17325 12328
rect 17359 12325 17371 12359
rect 17313 12319 17371 12325
rect 17034 12288 17040 12300
rect 16995 12260 17040 12288
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1578 7392 1584 7404
rect 1539 7364 1584 7392
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 1765 6987 1823 6993
rect 1765 6984 1777 6987
rect 1636 6956 1777 6984
rect 1636 6944 1642 6956
rect 1765 6953 1777 6956
rect 1811 6953 1823 6987
rect 1765 6947 1823 6953
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 37369 5831 37427 5837
rect 37369 5797 37381 5831
rect 37415 5797 37427 5831
rect 37369 5791 37427 5797
rect 37384 5760 37412 5791
rect 37384 5732 38056 5760
rect 37550 5692 37556 5704
rect 37511 5664 37556 5692
rect 37550 5652 37556 5664
rect 37608 5652 37614 5704
rect 38028 5701 38056 5732
rect 38013 5695 38071 5701
rect 38013 5661 38025 5695
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 38194 5556 38200 5568
rect 38155 5528 38200 5556
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 9122 3068 9128 3120
rect 9180 3108 9186 3120
rect 9180 3080 26234 3108
rect 9180 3068 9186 3080
rect 25593 3043 25651 3049
rect 25593 3009 25605 3043
rect 25639 3009 25651 3043
rect 26206 3040 26234 3080
rect 32493 3043 32551 3049
rect 32493 3040 32505 3043
rect 26206 3012 32505 3040
rect 25593 3003 25651 3009
rect 32493 3009 32505 3012
rect 32539 3040 32551 3043
rect 32769 3043 32827 3049
rect 32769 3040 32781 3043
rect 32539 3012 32781 3040
rect 32539 3009 32551 3012
rect 32493 3003 32551 3009
rect 32769 3009 32781 3012
rect 32815 3009 32827 3043
rect 32769 3003 32827 3009
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 25225 2907 25283 2913
rect 25225 2904 25237 2907
rect 9088 2876 25237 2904
rect 9088 2864 9094 2876
rect 25225 2873 25237 2876
rect 25271 2904 25283 2907
rect 25608 2904 25636 3003
rect 37550 2904 37556 2916
rect 25271 2876 37556 2904
rect 25271 2873 25283 2876
rect 25225 2867 25283 2873
rect 37550 2864 37556 2876
rect 37608 2864 37614 2916
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 25866 2836 25872 2848
rect 25823 2808 25872 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 32306 2836 32312 2848
rect 32267 2808 32312 2836
rect 32306 2796 32312 2808
rect 32364 2796 32370 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 6546 2632 6552 2644
rect 6507 2604 6552 2632
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 19429 2635 19487 2641
rect 19429 2632 19441 2635
rect 19392 2604 19441 2632
rect 19392 2592 19398 2604
rect 19429 2601 19441 2604
rect 19475 2601 19487 2635
rect 19429 2595 19487 2601
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 15286 2496 15292 2508
rect 1903 2468 15292 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 19426 2496 19432 2508
rect 16546 2468 19432 2496
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 72 2400 1593 2428
rect 72 2388 78 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6512 2400 6745 2428
rect 6512 2388 6518 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2428 13047 2431
rect 16546 2428 16574 2468
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 24820 2468 35894 2496
rect 24820 2456 24826 2468
rect 13035 2400 16574 2428
rect 13035 2397 13047 2400
rect 12989 2391 13047 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 25866 2428 25872 2440
rect 25827 2400 25872 2428
rect 19613 2391 19671 2397
rect 25866 2388 25872 2400
rect 25924 2388 25930 2440
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 35866 2428 35894 2468
rect 38013 2431 38071 2437
rect 38013 2428 38025 2431
rect 35866 2400 38025 2428
rect 38013 2397 38025 2400
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 32214 2252 32220 2304
rect 32272 2292 32278 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 32272 2264 32505 2292
rect 32272 2252 32278 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 38197 2295 38255 2301
rect 38197 2261 38209 2295
rect 38243 2292 38255 2295
rect 38654 2292 38660 2304
rect 38243 2264 38660 2292
rect 38243 2261 38255 2264
rect 38197 2255 38255 2261
rect 38654 2252 38660 2264
rect 38712 2252 38718 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 7104 37272 7156 37324
rect 664 37204 716 37256
rect 19432 37204 19484 37256
rect 19984 37204 20036 37256
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 32956 37247 33008 37256
rect 32956 37213 32965 37247
rect 32965 37213 32999 37247
rect 32999 37213 33008 37247
rect 32956 37204 33008 37213
rect 37832 37204 37884 37256
rect 7104 37136 7156 37188
rect 3792 37068 3844 37120
rect 13820 37068 13872 37120
rect 20076 37111 20128 37120
rect 20076 37077 20085 37111
rect 20085 37077 20119 37111
rect 20119 37077 20128 37111
rect 20076 37068 20128 37077
rect 26424 37068 26476 37120
rect 32864 37068 32916 37120
rect 39304 37068 39356 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 19432 36907 19484 36916
rect 19432 36873 19441 36907
rect 19441 36873 19475 36907
rect 19475 36873 19484 36907
rect 19432 36864 19484 36873
rect 20076 36728 20128 36780
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1676 34552 1728 34604
rect 1768 34391 1820 34400
rect 1768 34357 1777 34391
rect 1777 34357 1811 34391
rect 1811 34357 1820 34391
rect 1768 34348 1820 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 9864 33983 9916 33992
rect 9864 33949 9873 33983
rect 9873 33949 9907 33983
rect 9907 33949 9916 33983
rect 9864 33940 9916 33949
rect 12624 33940 12676 33992
rect 17316 34076 17368 34128
rect 13912 34008 13964 34060
rect 16212 34008 16264 34060
rect 14372 33983 14424 33992
rect 14372 33949 14381 33983
rect 14381 33949 14415 33983
rect 14415 33949 14424 33983
rect 14372 33940 14424 33949
rect 15476 33940 15528 33992
rect 15936 33983 15988 33992
rect 15936 33949 15945 33983
rect 15945 33949 15979 33983
rect 15979 33949 15988 33983
rect 15936 33940 15988 33949
rect 12900 33872 12952 33924
rect 9680 33847 9732 33856
rect 9680 33813 9689 33847
rect 9689 33813 9723 33847
rect 9723 33813 9732 33847
rect 9680 33804 9732 33813
rect 14004 33804 14056 33856
rect 14648 33847 14700 33856
rect 14648 33813 14657 33847
rect 14657 33813 14691 33847
rect 14691 33813 14700 33847
rect 14648 33804 14700 33813
rect 16120 33804 16172 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 15936 33600 15988 33652
rect 9680 33532 9732 33584
rect 8300 33464 8352 33516
rect 12624 33507 12676 33516
rect 12624 33473 12633 33507
rect 12633 33473 12667 33507
rect 12667 33473 12676 33507
rect 12624 33464 12676 33473
rect 13820 33464 13872 33516
rect 15292 33464 15344 33516
rect 8116 33260 8168 33312
rect 12072 33396 12124 33448
rect 14004 33439 14056 33448
rect 14004 33405 14013 33439
rect 14013 33405 14047 33439
rect 14047 33405 14056 33439
rect 14004 33396 14056 33405
rect 16212 33396 16264 33448
rect 8852 33303 8904 33312
rect 8852 33269 8861 33303
rect 8861 33269 8895 33303
rect 8895 33269 8904 33303
rect 8852 33260 8904 33269
rect 10968 33303 11020 33312
rect 10968 33269 10977 33303
rect 10977 33269 11011 33303
rect 11011 33269 11020 33303
rect 10968 33260 11020 33269
rect 12808 33260 12860 33312
rect 13912 33260 13964 33312
rect 17040 33328 17092 33380
rect 14924 33260 14976 33312
rect 15752 33260 15804 33312
rect 16488 33260 16540 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 9864 33056 9916 33108
rect 12808 33056 12860 33108
rect 12900 33056 12952 33108
rect 8852 32920 8904 32972
rect 15568 32963 15620 32972
rect 7472 32895 7524 32904
rect 7472 32861 7481 32895
rect 7481 32861 7515 32895
rect 7515 32861 7524 32895
rect 7472 32852 7524 32861
rect 8392 32895 8444 32904
rect 8392 32861 8401 32895
rect 8401 32861 8435 32895
rect 8435 32861 8444 32895
rect 8392 32852 8444 32861
rect 9404 32895 9456 32904
rect 9404 32861 9413 32895
rect 9413 32861 9447 32895
rect 9447 32861 9456 32895
rect 9404 32852 9456 32861
rect 10968 32852 11020 32904
rect 11060 32852 11112 32904
rect 12900 32852 12952 32904
rect 12716 32784 12768 32836
rect 7656 32759 7708 32768
rect 7656 32725 7665 32759
rect 7665 32725 7699 32759
rect 7699 32725 7708 32759
rect 7656 32716 7708 32725
rect 10324 32716 10376 32768
rect 14372 32852 14424 32904
rect 15568 32929 15577 32963
rect 15577 32929 15611 32963
rect 15611 32929 15620 32963
rect 15568 32920 15620 32929
rect 16672 33056 16724 33108
rect 15476 32852 15528 32904
rect 16120 32852 16172 32904
rect 38292 32895 38344 32904
rect 38292 32861 38301 32895
rect 38301 32861 38335 32895
rect 38335 32861 38344 32895
rect 38292 32852 38344 32861
rect 15384 32827 15436 32836
rect 15384 32793 15393 32827
rect 15393 32793 15427 32827
rect 15427 32793 15436 32827
rect 15384 32784 15436 32793
rect 18052 32784 18104 32836
rect 13544 32759 13596 32768
rect 13544 32725 13553 32759
rect 13553 32725 13587 32759
rect 13587 32725 13596 32759
rect 13544 32716 13596 32725
rect 14832 32759 14884 32768
rect 14832 32725 14841 32759
rect 14841 32725 14875 32759
rect 14875 32725 14884 32759
rect 14832 32716 14884 32725
rect 15476 32716 15528 32768
rect 16028 32716 16080 32768
rect 16764 32716 16816 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 7288 32512 7340 32564
rect 8116 32444 8168 32496
rect 8300 32512 8352 32564
rect 8760 32512 8812 32564
rect 11060 32512 11112 32564
rect 12716 32555 12768 32564
rect 12716 32521 12725 32555
rect 12725 32521 12759 32555
rect 12759 32521 12768 32555
rect 12716 32512 12768 32521
rect 14372 32512 14424 32564
rect 16028 32512 16080 32564
rect 6828 32419 6880 32428
rect 6828 32385 6862 32419
rect 6862 32385 6880 32419
rect 6828 32376 6880 32385
rect 7656 32376 7708 32428
rect 10324 32444 10376 32496
rect 9496 32376 9548 32428
rect 11060 32419 11112 32428
rect 8852 32308 8904 32360
rect 11060 32385 11069 32419
rect 11069 32385 11103 32419
rect 11103 32385 11112 32419
rect 11060 32376 11112 32385
rect 12716 32376 12768 32428
rect 13176 32376 13228 32428
rect 8576 32240 8628 32292
rect 9772 32283 9824 32292
rect 9772 32249 9781 32283
rect 9781 32249 9815 32283
rect 9815 32249 9824 32283
rect 9772 32240 9824 32249
rect 10968 32308 11020 32360
rect 11888 32240 11940 32292
rect 7932 32215 7984 32224
rect 7932 32181 7941 32215
rect 7941 32181 7975 32215
rect 7975 32181 7984 32215
rect 7932 32172 7984 32181
rect 10600 32172 10652 32224
rect 10968 32215 11020 32224
rect 10968 32181 10977 32215
rect 10977 32181 11011 32215
rect 11011 32181 11020 32215
rect 10968 32172 11020 32181
rect 11980 32172 12032 32224
rect 14648 32444 14700 32496
rect 15568 32444 15620 32496
rect 15476 32376 15528 32428
rect 15660 32419 15712 32428
rect 15660 32385 15669 32419
rect 15669 32385 15703 32419
rect 15703 32385 15712 32419
rect 15660 32376 15712 32385
rect 15844 32419 15896 32428
rect 15844 32385 15853 32419
rect 15853 32385 15887 32419
rect 15887 32385 15896 32419
rect 15844 32376 15896 32385
rect 16488 32376 16540 32428
rect 17224 32376 17276 32428
rect 13820 32240 13872 32292
rect 14556 32308 14608 32360
rect 15292 32308 15344 32360
rect 16764 32240 16816 32292
rect 14556 32172 14608 32224
rect 16212 32172 16264 32224
rect 17684 32215 17736 32224
rect 17684 32181 17693 32215
rect 17693 32181 17727 32215
rect 17727 32181 17736 32215
rect 17684 32172 17736 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 8668 31968 8720 32020
rect 9404 31968 9456 32020
rect 12992 32011 13044 32020
rect 6368 31900 6420 31952
rect 6460 31900 6512 31952
rect 7932 31900 7984 31952
rect 8576 31943 8628 31952
rect 8576 31909 8585 31943
rect 8585 31909 8619 31943
rect 8619 31909 8628 31943
rect 8576 31900 8628 31909
rect 9220 31900 9272 31952
rect 12992 31977 13001 32011
rect 13001 31977 13035 32011
rect 13035 31977 13044 32011
rect 12992 31968 13044 31977
rect 13176 32011 13228 32020
rect 13176 31977 13185 32011
rect 13185 31977 13219 32011
rect 13219 31977 13228 32011
rect 13176 31968 13228 31977
rect 27160 31968 27212 32020
rect 14372 31900 14424 31952
rect 2780 31764 2832 31816
rect 5172 31807 5224 31816
rect 2504 31696 2556 31748
rect 5172 31773 5181 31807
rect 5181 31773 5215 31807
rect 5215 31773 5224 31807
rect 5172 31764 5224 31773
rect 9680 31832 9732 31884
rect 10324 31875 10376 31884
rect 10324 31841 10333 31875
rect 10333 31841 10367 31875
rect 10367 31841 10376 31875
rect 10324 31832 10376 31841
rect 10968 31832 11020 31884
rect 11888 31875 11940 31884
rect 5816 31807 5868 31816
rect 5816 31773 5825 31807
rect 5825 31773 5859 31807
rect 5859 31773 5868 31807
rect 5816 31764 5868 31773
rect 6460 31807 6512 31816
rect 5448 31696 5500 31748
rect 6460 31773 6469 31807
rect 6469 31773 6503 31807
rect 6503 31773 6512 31807
rect 6460 31764 6512 31773
rect 6644 31764 6696 31816
rect 8024 31764 8076 31816
rect 9588 31764 9640 31816
rect 10140 31764 10192 31816
rect 10600 31807 10652 31816
rect 10600 31773 10609 31807
rect 10609 31773 10643 31807
rect 10643 31773 10652 31807
rect 10600 31764 10652 31773
rect 11060 31764 11112 31816
rect 11152 31764 11204 31816
rect 11888 31841 11897 31875
rect 11897 31841 11931 31875
rect 11931 31841 11940 31875
rect 11888 31832 11940 31841
rect 12716 31832 12768 31884
rect 14188 31832 14240 31884
rect 15476 31875 15528 31884
rect 14372 31764 14424 31816
rect 14648 31807 14700 31816
rect 14648 31773 14657 31807
rect 14657 31773 14691 31807
rect 14691 31773 14700 31807
rect 14648 31764 14700 31773
rect 15476 31841 15485 31875
rect 15485 31841 15519 31875
rect 15519 31841 15528 31875
rect 15476 31832 15528 31841
rect 15936 31900 15988 31952
rect 18052 31943 18104 31952
rect 18052 31909 18061 31943
rect 18061 31909 18095 31943
rect 18095 31909 18104 31943
rect 18052 31900 18104 31909
rect 15660 31875 15712 31884
rect 15660 31841 15669 31875
rect 15669 31841 15703 31875
rect 15703 31841 15712 31875
rect 15660 31832 15712 31841
rect 15844 31832 15896 31884
rect 17684 31764 17736 31816
rect 19984 31807 20036 31816
rect 19984 31773 19993 31807
rect 19993 31773 20027 31807
rect 20027 31773 20036 31807
rect 19984 31764 20036 31773
rect 8300 31696 8352 31748
rect 5908 31671 5960 31680
rect 5908 31637 5917 31671
rect 5917 31637 5951 31671
rect 5951 31637 5960 31671
rect 5908 31628 5960 31637
rect 6000 31628 6052 31680
rect 11244 31696 11296 31748
rect 11980 31739 12032 31748
rect 11980 31705 11989 31739
rect 11989 31705 12023 31739
rect 12023 31705 12032 31739
rect 11980 31696 12032 31705
rect 13728 31696 13780 31748
rect 14464 31739 14516 31748
rect 14464 31705 14473 31739
rect 14473 31705 14507 31739
rect 14507 31705 14516 31739
rect 14464 31696 14516 31705
rect 14556 31739 14608 31748
rect 14556 31705 14565 31739
rect 14565 31705 14599 31739
rect 14599 31705 14608 31739
rect 14556 31696 14608 31705
rect 15476 31696 15528 31748
rect 9956 31628 10008 31680
rect 10692 31671 10744 31680
rect 10692 31637 10701 31671
rect 10701 31637 10735 31671
rect 10735 31637 10744 31671
rect 10692 31628 10744 31637
rect 11336 31671 11388 31680
rect 11336 31637 11345 31671
rect 11345 31637 11379 31671
rect 11379 31637 11388 31671
rect 11336 31628 11388 31637
rect 11520 31628 11572 31680
rect 12440 31628 12492 31680
rect 15292 31671 15344 31680
rect 15292 31637 15301 31671
rect 15301 31637 15335 31671
rect 15335 31637 15344 31671
rect 15292 31628 15344 31637
rect 20076 31628 20128 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1952 31220 2004 31272
rect 2504 31263 2556 31272
rect 2504 31229 2513 31263
rect 2513 31229 2547 31263
rect 2547 31229 2556 31263
rect 2504 31220 2556 31229
rect 2596 31220 2648 31272
rect 2780 31356 2832 31408
rect 5816 31424 5868 31476
rect 6736 31467 6788 31476
rect 6736 31433 6745 31467
rect 6745 31433 6779 31467
rect 6779 31433 6788 31467
rect 6736 31424 6788 31433
rect 8116 31424 8168 31476
rect 3792 31331 3844 31340
rect 3792 31297 3801 31331
rect 3801 31297 3835 31331
rect 3835 31297 3844 31331
rect 3792 31288 3844 31297
rect 4988 31288 5040 31340
rect 6000 31288 6052 31340
rect 6644 31331 6696 31340
rect 6644 31297 6653 31331
rect 6653 31297 6687 31331
rect 6687 31297 6696 31331
rect 6644 31288 6696 31297
rect 7288 31331 7340 31340
rect 6460 31220 6512 31272
rect 7288 31297 7297 31331
rect 7297 31297 7331 31331
rect 7331 31297 7340 31331
rect 7288 31288 7340 31297
rect 8024 31288 8076 31340
rect 8297 31331 8349 31340
rect 8297 31297 8306 31331
rect 8306 31297 8340 31331
rect 8340 31297 8349 31331
rect 8297 31288 8349 31297
rect 8668 31288 8720 31340
rect 9772 31356 9824 31408
rect 10784 31399 10836 31408
rect 10784 31365 10793 31399
rect 10793 31365 10827 31399
rect 10827 31365 10836 31399
rect 10784 31356 10836 31365
rect 10968 31399 11020 31408
rect 10968 31365 11003 31399
rect 11003 31365 11020 31399
rect 10968 31356 11020 31365
rect 11244 31356 11296 31408
rect 12164 31356 12216 31408
rect 9680 31331 9732 31340
rect 9680 31297 9689 31331
rect 9689 31297 9723 31331
rect 9723 31297 9732 31331
rect 9680 31288 9732 31297
rect 9864 31331 9916 31340
rect 9864 31297 9873 31331
rect 9873 31297 9907 31331
rect 9907 31297 9916 31331
rect 9864 31288 9916 31297
rect 10600 31288 10652 31340
rect 11888 31331 11940 31340
rect 11888 31297 11897 31331
rect 11897 31297 11931 31331
rect 11931 31297 11940 31331
rect 11888 31288 11940 31297
rect 12440 31467 12492 31476
rect 12440 31433 12449 31467
rect 12449 31433 12483 31467
rect 12483 31433 12492 31467
rect 12440 31424 12492 31433
rect 13268 31399 13320 31408
rect 13268 31365 13277 31399
rect 13277 31365 13311 31399
rect 13311 31365 13320 31399
rect 13268 31356 13320 31365
rect 20076 31399 20128 31408
rect 20076 31365 20110 31399
rect 20110 31365 20128 31399
rect 20076 31356 20128 31365
rect 25320 31356 25372 31408
rect 13084 31331 13136 31340
rect 13084 31297 13093 31331
rect 13093 31297 13127 31331
rect 13127 31297 13136 31331
rect 13084 31288 13136 31297
rect 13176 31331 13228 31340
rect 13176 31297 13185 31331
rect 13185 31297 13219 31331
rect 13219 31297 13228 31331
rect 13176 31288 13228 31297
rect 14372 31288 14424 31340
rect 16304 31331 16356 31340
rect 16304 31297 16313 31331
rect 16313 31297 16347 31331
rect 16347 31297 16356 31331
rect 16304 31288 16356 31297
rect 17316 31331 17368 31340
rect 17316 31297 17325 31331
rect 17325 31297 17359 31331
rect 17359 31297 17368 31331
rect 17316 31288 17368 31297
rect 17868 31288 17920 31340
rect 22008 31331 22060 31340
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 23112 31331 23164 31340
rect 23112 31297 23121 31331
rect 23121 31297 23155 31331
rect 23155 31297 23164 31331
rect 23112 31288 23164 31297
rect 23388 31331 23440 31340
rect 23388 31297 23397 31331
rect 23397 31297 23431 31331
rect 23431 31297 23440 31331
rect 23388 31288 23440 31297
rect 8760 31220 8812 31272
rect 9496 31220 9548 31272
rect 11152 31263 11204 31272
rect 11152 31229 11161 31263
rect 11161 31229 11195 31263
rect 11195 31229 11204 31263
rect 11152 31220 11204 31229
rect 11244 31220 11296 31272
rect 6552 31152 6604 31204
rect 8576 31152 8628 31204
rect 5724 31084 5776 31136
rect 7748 31084 7800 31136
rect 8024 31084 8076 31136
rect 10048 31127 10100 31136
rect 10048 31093 10057 31127
rect 10057 31093 10091 31127
rect 10091 31093 10100 31127
rect 10048 31084 10100 31093
rect 11336 31084 11388 31136
rect 13544 31152 13596 31204
rect 14372 31152 14424 31204
rect 18972 31220 19024 31272
rect 24860 31288 24912 31340
rect 24768 31263 24820 31272
rect 24768 31229 24777 31263
rect 24777 31229 24811 31263
rect 24811 31229 24820 31263
rect 24768 31220 24820 31229
rect 14464 31084 14516 31136
rect 14832 31084 14884 31136
rect 16028 31084 16080 31136
rect 16948 31084 17000 31136
rect 18880 31084 18932 31136
rect 19432 31084 19484 31136
rect 23020 31152 23072 31204
rect 32956 31152 33008 31204
rect 20904 31084 20956 31136
rect 22008 31084 22060 31136
rect 22284 31127 22336 31136
rect 22284 31093 22293 31127
rect 22293 31093 22327 31127
rect 22327 31093 22336 31127
rect 22284 31084 22336 31093
rect 23204 31084 23256 31136
rect 24676 31127 24728 31136
rect 24676 31093 24685 31127
rect 24685 31093 24719 31127
rect 24719 31093 24728 31127
rect 24676 31084 24728 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2596 30744 2648 30796
rect 2136 30676 2188 30728
rect 5724 30744 5776 30796
rect 6644 30812 6696 30864
rect 11704 30880 11756 30932
rect 11888 30923 11940 30932
rect 11888 30889 11897 30923
rect 11897 30889 11931 30923
rect 11931 30889 11940 30923
rect 11888 30880 11940 30889
rect 12992 30880 13044 30932
rect 15292 30880 15344 30932
rect 10048 30812 10100 30864
rect 15752 30880 15804 30932
rect 16212 30880 16264 30932
rect 17224 30880 17276 30932
rect 17868 30923 17920 30932
rect 17868 30889 17877 30923
rect 17877 30889 17911 30923
rect 17911 30889 17920 30923
rect 17868 30880 17920 30889
rect 24676 30880 24728 30932
rect 4804 30719 4856 30728
rect 4804 30685 4813 30719
rect 4813 30685 4847 30719
rect 4847 30685 4856 30719
rect 4804 30676 4856 30685
rect 5448 30676 5500 30728
rect 6736 30744 6788 30796
rect 7748 30719 7800 30728
rect 7748 30685 7757 30719
rect 7757 30685 7791 30719
rect 7791 30685 7800 30719
rect 7748 30676 7800 30685
rect 8300 30744 8352 30796
rect 8484 30744 8536 30796
rect 9496 30744 9548 30796
rect 8024 30719 8076 30728
rect 8024 30685 8033 30719
rect 8033 30685 8067 30719
rect 8067 30685 8076 30719
rect 8024 30676 8076 30685
rect 7380 30608 7432 30660
rect 4436 30583 4488 30592
rect 4436 30549 4445 30583
rect 4445 30549 4479 30583
rect 4479 30549 4488 30583
rect 4436 30540 4488 30549
rect 5816 30540 5868 30592
rect 8576 30540 8628 30592
rect 9588 30719 9640 30728
rect 9588 30685 9597 30719
rect 9597 30685 9631 30719
rect 9631 30685 9640 30719
rect 9588 30676 9640 30685
rect 9956 30744 10008 30796
rect 10600 30787 10652 30796
rect 10140 30676 10192 30728
rect 10324 30719 10376 30728
rect 10324 30685 10333 30719
rect 10333 30685 10367 30719
rect 10367 30685 10376 30719
rect 10324 30676 10376 30685
rect 10600 30753 10609 30787
rect 10609 30753 10643 30787
rect 10643 30753 10652 30787
rect 10600 30744 10652 30753
rect 15844 30812 15896 30864
rect 19984 30812 20036 30864
rect 11428 30787 11480 30796
rect 11428 30753 11437 30787
rect 11437 30753 11471 30787
rect 11471 30753 11480 30787
rect 11428 30744 11480 30753
rect 11612 30744 11664 30796
rect 12716 30787 12768 30796
rect 12716 30753 12725 30787
rect 12725 30753 12759 30787
rect 12759 30753 12768 30787
rect 12716 30744 12768 30753
rect 13452 30744 13504 30796
rect 14372 30744 14424 30796
rect 20904 30787 20956 30796
rect 20904 30753 20913 30787
rect 20913 30753 20947 30787
rect 20947 30753 20956 30787
rect 20904 30744 20956 30753
rect 21180 30787 21232 30796
rect 9864 30608 9916 30660
rect 9772 30540 9824 30592
rect 10600 30540 10652 30592
rect 11060 30540 11112 30592
rect 11520 30719 11572 30728
rect 11520 30685 11529 30719
rect 11529 30685 11563 30719
rect 11563 30685 11572 30719
rect 11520 30676 11572 30685
rect 11796 30676 11848 30728
rect 12992 30676 13044 30728
rect 13176 30719 13228 30728
rect 13176 30685 13185 30719
rect 13185 30685 13219 30719
rect 13219 30685 13228 30719
rect 13176 30676 13228 30685
rect 16028 30676 16080 30728
rect 17040 30719 17092 30728
rect 13728 30608 13780 30660
rect 13084 30583 13136 30592
rect 13084 30549 13093 30583
rect 13093 30549 13127 30583
rect 13127 30549 13136 30583
rect 13084 30540 13136 30549
rect 14648 30583 14700 30592
rect 14648 30549 14673 30583
rect 14673 30549 14700 30583
rect 14832 30583 14884 30592
rect 14648 30540 14700 30549
rect 14832 30549 14841 30583
rect 14841 30549 14875 30583
rect 14875 30549 14884 30583
rect 14832 30540 14884 30549
rect 15292 30651 15344 30660
rect 15292 30617 15301 30651
rect 15301 30617 15335 30651
rect 15335 30617 15344 30651
rect 15292 30608 15344 30617
rect 15651 30608 15703 30660
rect 17040 30685 17049 30719
rect 17049 30685 17083 30719
rect 17083 30685 17092 30719
rect 17040 30676 17092 30685
rect 18420 30676 18472 30728
rect 20444 30719 20496 30728
rect 20444 30685 20453 30719
rect 20453 30685 20487 30719
rect 20487 30685 20496 30719
rect 20444 30676 20496 30685
rect 19248 30608 19300 30660
rect 19340 30608 19392 30660
rect 21180 30753 21189 30787
rect 21189 30753 21223 30787
rect 21223 30753 21232 30787
rect 21180 30744 21232 30753
rect 23020 30787 23072 30796
rect 23020 30753 23029 30787
rect 23029 30753 23063 30787
rect 23063 30753 23072 30787
rect 23020 30744 23072 30753
rect 22560 30676 22612 30728
rect 24676 30676 24728 30728
rect 25044 30719 25096 30728
rect 25044 30685 25053 30719
rect 25053 30685 25087 30719
rect 25087 30685 25096 30719
rect 25044 30676 25096 30685
rect 18696 30583 18748 30592
rect 18696 30549 18721 30583
rect 18721 30549 18748 30583
rect 18696 30540 18748 30549
rect 19064 30540 19116 30592
rect 20352 30540 20404 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4436 30379 4488 30388
rect 4436 30345 4445 30379
rect 4445 30345 4479 30379
rect 4479 30345 4488 30379
rect 4436 30336 4488 30345
rect 5816 30379 5868 30388
rect 5816 30345 5825 30379
rect 5825 30345 5859 30379
rect 5859 30345 5868 30379
rect 5816 30336 5868 30345
rect 6552 30336 6604 30388
rect 8484 30379 8536 30388
rect 4620 30268 4672 30320
rect 6828 30311 6880 30320
rect 6828 30277 6837 30311
rect 6837 30277 6871 30311
rect 6871 30277 6880 30311
rect 6828 30268 6880 30277
rect 8484 30345 8493 30379
rect 8493 30345 8527 30379
rect 8527 30345 8536 30379
rect 8484 30336 8536 30345
rect 9956 30336 10008 30388
rect 10692 30336 10744 30388
rect 13176 30336 13228 30388
rect 16304 30379 16356 30388
rect 16304 30345 16313 30379
rect 16313 30345 16347 30379
rect 16347 30345 16356 30379
rect 16304 30336 16356 30345
rect 18696 30336 18748 30388
rect 23112 30336 23164 30388
rect 24676 30336 24728 30388
rect 2688 30243 2740 30252
rect 2688 30209 2722 30243
rect 2722 30209 2740 30243
rect 2688 30200 2740 30209
rect 4068 30200 4120 30252
rect 2136 30132 2188 30184
rect 6368 30200 6420 30252
rect 6644 30243 6696 30252
rect 6644 30209 6653 30243
rect 6653 30209 6687 30243
rect 6687 30209 6696 30243
rect 7564 30311 7616 30320
rect 7564 30277 7573 30311
rect 7573 30277 7607 30311
rect 7607 30277 7616 30311
rect 7564 30268 7616 30277
rect 9404 30268 9456 30320
rect 11520 30268 11572 30320
rect 14188 30311 14240 30320
rect 14188 30277 14197 30311
rect 14197 30277 14231 30311
rect 14231 30277 14240 30311
rect 14188 30268 14240 30277
rect 14556 30311 14608 30320
rect 14556 30277 14565 30311
rect 14565 30277 14599 30311
rect 14599 30277 14608 30311
rect 14556 30268 14608 30277
rect 16028 30268 16080 30320
rect 17316 30268 17368 30320
rect 22008 30311 22060 30320
rect 6644 30200 6696 30209
rect 9220 30243 9272 30252
rect 6736 30132 6788 30184
rect 6828 30175 6880 30184
rect 6828 30141 6837 30175
rect 6837 30141 6871 30175
rect 6871 30141 6880 30175
rect 6828 30132 6880 30141
rect 8024 30132 8076 30184
rect 9220 30209 9229 30243
rect 9229 30209 9263 30243
rect 9263 30209 9272 30243
rect 9220 30200 9272 30209
rect 7564 30064 7616 30116
rect 11612 30200 11664 30252
rect 10600 30132 10652 30184
rect 13544 30243 13596 30252
rect 13544 30209 13553 30243
rect 13553 30209 13587 30243
rect 13587 30209 13596 30243
rect 13544 30200 13596 30209
rect 12256 30175 12308 30184
rect 12256 30141 12265 30175
rect 12265 30141 12299 30175
rect 12299 30141 12308 30175
rect 12256 30132 12308 30141
rect 12532 30175 12584 30184
rect 12532 30141 12541 30175
rect 12541 30141 12575 30175
rect 12575 30141 12584 30175
rect 12532 30132 12584 30141
rect 12992 30132 13044 30184
rect 13636 30132 13688 30184
rect 3884 29996 3936 30048
rect 5172 29996 5224 30048
rect 5816 29996 5868 30048
rect 6644 29996 6696 30048
rect 6828 29996 6880 30048
rect 7932 29996 7984 30048
rect 13544 30064 13596 30116
rect 14464 30243 14516 30252
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 15752 30243 15804 30252
rect 14464 30200 14516 30209
rect 15752 30209 15761 30243
rect 15761 30209 15795 30243
rect 15795 30209 15804 30243
rect 15752 30200 15804 30209
rect 16672 30200 16724 30252
rect 16948 30200 17000 30252
rect 19064 30243 19116 30252
rect 15108 30132 15160 30184
rect 15568 30132 15620 30184
rect 19064 30209 19073 30243
rect 19073 30209 19107 30243
rect 19107 30209 19116 30243
rect 19064 30200 19116 30209
rect 22008 30277 22017 30311
rect 22017 30277 22051 30311
rect 22051 30277 22060 30311
rect 22008 30268 22060 30277
rect 25320 30311 25372 30320
rect 25320 30277 25329 30311
rect 25329 30277 25363 30311
rect 25363 30277 25372 30311
rect 25320 30268 25372 30277
rect 20352 30243 20404 30252
rect 20352 30209 20386 30243
rect 20386 30209 20404 30243
rect 20352 30200 20404 30209
rect 22560 30200 22612 30252
rect 19340 30132 19392 30184
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 24584 30132 24636 30184
rect 25044 30175 25096 30184
rect 25044 30141 25053 30175
rect 25053 30141 25087 30175
rect 25087 30141 25096 30175
rect 25044 30132 25096 30141
rect 15844 30064 15896 30116
rect 22284 30107 22336 30116
rect 22284 30073 22293 30107
rect 22293 30073 22327 30107
rect 22327 30073 22336 30107
rect 22284 30064 22336 30073
rect 10968 29996 11020 30048
rect 12624 29996 12676 30048
rect 14464 29996 14516 30048
rect 15292 29996 15344 30048
rect 15752 29996 15804 30048
rect 16488 29996 16540 30048
rect 17132 29996 17184 30048
rect 21456 30039 21508 30048
rect 21456 30005 21465 30039
rect 21465 30005 21499 30039
rect 21499 30005 21508 30039
rect 21456 29996 21508 30005
rect 25044 29996 25096 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2688 29792 2740 29844
rect 4068 29792 4120 29844
rect 4160 29792 4212 29844
rect 8024 29792 8076 29844
rect 11244 29792 11296 29844
rect 12072 29792 12124 29844
rect 3884 29656 3936 29708
rect 2688 29588 2740 29640
rect 9220 29724 9272 29776
rect 14372 29792 14424 29844
rect 14648 29792 14700 29844
rect 15016 29792 15068 29844
rect 15476 29835 15528 29844
rect 15476 29801 15485 29835
rect 15485 29801 15519 29835
rect 15519 29801 15528 29835
rect 15476 29792 15528 29801
rect 16028 29835 16080 29844
rect 16028 29801 16037 29835
rect 16037 29801 16071 29835
rect 16071 29801 16080 29835
rect 16028 29792 16080 29801
rect 16488 29792 16540 29844
rect 18420 29835 18472 29844
rect 12532 29767 12584 29776
rect 12532 29733 12541 29767
rect 12541 29733 12575 29767
rect 12575 29733 12584 29767
rect 12532 29724 12584 29733
rect 4620 29656 4672 29708
rect 5448 29656 5500 29708
rect 5908 29656 5960 29708
rect 8116 29656 8168 29708
rect 10324 29656 10376 29708
rect 10508 29656 10560 29708
rect 12072 29699 12124 29708
rect 5356 29588 5408 29640
rect 5540 29631 5592 29640
rect 5540 29597 5549 29631
rect 5549 29597 5583 29631
rect 5583 29597 5592 29631
rect 5540 29588 5592 29597
rect 4804 29520 4856 29572
rect 7288 29588 7340 29640
rect 8208 29631 8260 29640
rect 8208 29597 8217 29631
rect 8217 29597 8251 29631
rect 8251 29597 8260 29631
rect 8208 29588 8260 29597
rect 9128 29631 9180 29640
rect 9128 29597 9137 29631
rect 9137 29597 9171 29631
rect 9171 29597 9180 29631
rect 9128 29588 9180 29597
rect 9312 29631 9364 29640
rect 9312 29597 9340 29631
rect 9340 29597 9364 29631
rect 9312 29588 9364 29597
rect 9588 29588 9640 29640
rect 12072 29665 12081 29699
rect 12081 29665 12115 29699
rect 12115 29665 12124 29699
rect 12072 29656 12124 29665
rect 14740 29724 14792 29776
rect 15292 29724 15344 29776
rect 18420 29801 18429 29835
rect 18429 29801 18463 29835
rect 18463 29801 18472 29835
rect 18420 29792 18472 29801
rect 20444 29792 20496 29844
rect 21180 29835 21232 29844
rect 21180 29801 21189 29835
rect 21189 29801 21223 29835
rect 21223 29801 21232 29835
rect 21180 29792 21232 29801
rect 23388 29792 23440 29844
rect 24860 29792 24912 29844
rect 23296 29724 23348 29776
rect 6828 29563 6880 29572
rect 6828 29529 6837 29563
rect 6837 29529 6871 29563
rect 6871 29529 6880 29563
rect 6828 29520 6880 29529
rect 7012 29563 7064 29572
rect 7012 29529 7021 29563
rect 7021 29529 7055 29563
rect 7055 29529 7064 29563
rect 7012 29520 7064 29529
rect 8760 29520 8812 29572
rect 10784 29631 10836 29640
rect 10784 29597 10793 29631
rect 10793 29597 10827 29631
rect 10827 29597 10836 29631
rect 10784 29588 10836 29597
rect 10968 29631 11020 29640
rect 10968 29597 10977 29631
rect 10977 29597 11011 29631
rect 11011 29597 11020 29631
rect 13636 29656 13688 29708
rect 10968 29588 11020 29597
rect 11888 29520 11940 29572
rect 7196 29495 7248 29504
rect 7196 29461 7205 29495
rect 7205 29461 7239 29495
rect 7239 29461 7248 29495
rect 7196 29452 7248 29461
rect 8576 29495 8628 29504
rect 8576 29461 8585 29495
rect 8585 29461 8619 29495
rect 8619 29461 8628 29495
rect 8576 29452 8628 29461
rect 9496 29495 9548 29504
rect 9496 29461 9505 29495
rect 9505 29461 9539 29495
rect 9539 29461 9548 29495
rect 9496 29452 9548 29461
rect 10692 29452 10744 29504
rect 12348 29588 12400 29640
rect 13084 29588 13136 29640
rect 13728 29588 13780 29640
rect 19340 29656 19392 29708
rect 14556 29588 14608 29640
rect 14740 29588 14792 29640
rect 15292 29631 15344 29640
rect 15292 29597 15301 29631
rect 15301 29597 15335 29631
rect 15335 29597 15344 29631
rect 15292 29588 15344 29597
rect 15752 29588 15804 29640
rect 16488 29631 16540 29640
rect 16488 29597 16497 29631
rect 16497 29597 16531 29631
rect 16531 29597 16540 29631
rect 16488 29588 16540 29597
rect 15660 29520 15712 29572
rect 21456 29520 21508 29572
rect 23020 29588 23072 29640
rect 25044 29631 25096 29640
rect 25044 29597 25053 29631
rect 25053 29597 25087 29631
rect 25087 29597 25096 29631
rect 25044 29588 25096 29597
rect 25136 29520 25188 29572
rect 12532 29452 12584 29504
rect 14464 29495 14516 29504
rect 14464 29461 14473 29495
rect 14473 29461 14507 29495
rect 14507 29461 14516 29495
rect 14464 29452 14516 29461
rect 14556 29452 14608 29504
rect 16304 29452 16356 29504
rect 17868 29452 17920 29504
rect 20076 29452 20128 29504
rect 20536 29452 20588 29504
rect 21548 29452 21600 29504
rect 24676 29452 24728 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 7012 29248 7064 29300
rect 8392 29248 8444 29300
rect 10784 29248 10836 29300
rect 13268 29248 13320 29300
rect 8576 29180 8628 29232
rect 3516 29112 3568 29164
rect 6736 29155 6788 29164
rect 6736 29121 6745 29155
rect 6745 29121 6779 29155
rect 6779 29121 6788 29155
rect 6736 29112 6788 29121
rect 8300 29155 8352 29164
rect 4896 29044 4948 29096
rect 5356 29044 5408 29096
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 8300 29112 8352 29121
rect 8392 29155 8444 29164
rect 8392 29121 8401 29155
rect 8401 29121 8435 29155
rect 8435 29121 8444 29155
rect 9312 29180 9364 29232
rect 9496 29180 9548 29232
rect 12624 29223 12676 29232
rect 12624 29189 12633 29223
rect 12633 29189 12667 29223
rect 12667 29189 12676 29223
rect 12624 29180 12676 29189
rect 13544 29180 13596 29232
rect 15292 29248 15344 29300
rect 16212 29248 16264 29300
rect 17868 29291 17920 29300
rect 17868 29257 17877 29291
rect 17877 29257 17911 29291
rect 17911 29257 17920 29291
rect 17868 29248 17920 29257
rect 20076 29291 20128 29300
rect 15752 29180 15804 29232
rect 17592 29180 17644 29232
rect 8392 29112 8444 29121
rect 10324 29155 10376 29164
rect 10324 29121 10333 29155
rect 10333 29121 10367 29155
rect 10367 29121 10376 29155
rect 10324 29112 10376 29121
rect 11704 29155 11756 29164
rect 11704 29121 11713 29155
rect 11713 29121 11747 29155
rect 11747 29121 11756 29155
rect 11704 29112 11756 29121
rect 11888 29155 11940 29164
rect 11888 29121 11897 29155
rect 11897 29121 11931 29155
rect 11931 29121 11940 29155
rect 11888 29112 11940 29121
rect 12440 29112 12492 29164
rect 4160 29019 4212 29028
rect 4160 28985 4169 29019
rect 4169 28985 4203 29019
rect 4203 28985 4212 29019
rect 4160 28976 4212 28985
rect 8668 29044 8720 29096
rect 9128 29044 9180 29096
rect 8484 28976 8536 29028
rect 9496 29087 9548 29096
rect 9496 29053 9505 29087
rect 9505 29053 9539 29087
rect 9539 29053 9548 29087
rect 10600 29087 10652 29096
rect 9496 29044 9548 29053
rect 10600 29053 10609 29087
rect 10609 29053 10643 29087
rect 10643 29053 10652 29087
rect 10600 29044 10652 29053
rect 14740 29112 14792 29164
rect 14924 29155 14976 29164
rect 14924 29121 14933 29155
rect 14933 29121 14967 29155
rect 14967 29121 14976 29155
rect 14924 29112 14976 29121
rect 16764 29112 16816 29164
rect 17132 29112 17184 29164
rect 18236 29155 18288 29164
rect 18236 29121 18245 29155
rect 18245 29121 18279 29155
rect 18279 29121 18288 29155
rect 18236 29112 18288 29121
rect 17960 29044 18012 29096
rect 20076 29257 20085 29291
rect 20085 29257 20119 29291
rect 20119 29257 20128 29291
rect 20076 29248 20128 29257
rect 25044 29248 25096 29300
rect 19156 29180 19208 29232
rect 22744 29180 22796 29232
rect 20536 29155 20588 29164
rect 19432 29044 19484 29096
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 20904 29112 20956 29164
rect 21180 29155 21232 29164
rect 21180 29121 21189 29155
rect 21189 29121 21223 29155
rect 21223 29121 21232 29155
rect 21180 29112 21232 29121
rect 21456 29112 21508 29164
rect 22100 29112 22152 29164
rect 23112 29112 23164 29164
rect 22928 29087 22980 29096
rect 22928 29053 22937 29087
rect 22937 29053 22971 29087
rect 22971 29053 22980 29087
rect 22928 29044 22980 29053
rect 10968 28976 11020 29028
rect 12256 28976 12308 29028
rect 8300 28908 8352 28960
rect 9588 28908 9640 28960
rect 11888 28908 11940 28960
rect 19340 28976 19392 29028
rect 20536 28976 20588 29028
rect 25044 29044 25096 29096
rect 18236 28908 18288 28960
rect 20996 28951 21048 28960
rect 20996 28917 21005 28951
rect 21005 28917 21039 28951
rect 21039 28917 21048 28951
rect 20996 28908 21048 28917
rect 22376 28951 22428 28960
rect 22376 28917 22385 28951
rect 22385 28917 22419 28951
rect 22419 28917 22428 28951
rect 22376 28908 22428 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4896 28704 4948 28756
rect 4160 28543 4212 28552
rect 4160 28509 4169 28543
rect 4169 28509 4203 28543
rect 4203 28509 4212 28543
rect 4160 28500 4212 28509
rect 5264 28704 5316 28756
rect 5356 28500 5408 28552
rect 3976 28364 4028 28416
rect 5264 28364 5316 28416
rect 7472 28704 7524 28756
rect 6920 28636 6972 28688
rect 8392 28704 8444 28756
rect 8760 28704 8812 28756
rect 9404 28747 9456 28756
rect 9404 28713 9413 28747
rect 9413 28713 9447 28747
rect 9447 28713 9456 28747
rect 9404 28704 9456 28713
rect 9588 28747 9640 28756
rect 9588 28713 9597 28747
rect 9597 28713 9631 28747
rect 9631 28713 9640 28747
rect 9588 28704 9640 28713
rect 11888 28704 11940 28756
rect 14280 28704 14332 28756
rect 17040 28704 17092 28756
rect 25044 28747 25096 28756
rect 25044 28713 25053 28747
rect 25053 28713 25087 28747
rect 25087 28713 25096 28747
rect 25044 28704 25096 28713
rect 6828 28500 6880 28552
rect 7196 28568 7248 28620
rect 14648 28636 14700 28688
rect 18328 28636 18380 28688
rect 18788 28679 18840 28688
rect 18788 28645 18797 28679
rect 18797 28645 18831 28679
rect 18831 28645 18840 28679
rect 18788 28636 18840 28645
rect 19064 28636 19116 28688
rect 20904 28636 20956 28688
rect 7288 28500 7340 28552
rect 10508 28568 10560 28620
rect 8024 28543 8076 28552
rect 8024 28509 8033 28543
rect 8033 28509 8067 28543
rect 8067 28509 8076 28543
rect 8024 28500 8076 28509
rect 8484 28500 8536 28552
rect 9680 28500 9732 28552
rect 10600 28543 10652 28552
rect 10600 28509 10609 28543
rect 10609 28509 10643 28543
rect 10643 28509 10652 28543
rect 10600 28500 10652 28509
rect 10692 28500 10744 28552
rect 14740 28611 14792 28620
rect 14740 28577 14749 28611
rect 14749 28577 14783 28611
rect 14783 28577 14792 28611
rect 14740 28568 14792 28577
rect 14556 28543 14608 28552
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 6736 28432 6788 28484
rect 8760 28432 8812 28484
rect 12808 28432 12860 28484
rect 15016 28500 15068 28552
rect 15384 28500 15436 28552
rect 16580 28568 16632 28620
rect 16764 28568 16816 28620
rect 20720 28568 20772 28620
rect 15200 28475 15252 28484
rect 15200 28441 15209 28475
rect 15209 28441 15243 28475
rect 15243 28441 15252 28475
rect 15200 28432 15252 28441
rect 17960 28500 18012 28552
rect 18972 28500 19024 28552
rect 22928 28636 22980 28688
rect 23020 28611 23072 28620
rect 23020 28577 23029 28611
rect 23029 28577 23063 28611
rect 23063 28577 23072 28611
rect 23020 28568 23072 28577
rect 22192 28543 22244 28552
rect 18144 28432 18196 28484
rect 19432 28432 19484 28484
rect 11796 28364 11848 28416
rect 14648 28364 14700 28416
rect 15292 28407 15344 28416
rect 15292 28373 15301 28407
rect 15301 28373 15335 28407
rect 15335 28373 15344 28407
rect 15292 28364 15344 28373
rect 16396 28407 16448 28416
rect 16396 28373 16405 28407
rect 16405 28373 16439 28407
rect 16439 28373 16448 28407
rect 16396 28364 16448 28373
rect 17224 28364 17276 28416
rect 22192 28509 22201 28543
rect 22201 28509 22235 28543
rect 22235 28509 22244 28543
rect 22192 28500 22244 28509
rect 22376 28543 22428 28552
rect 22376 28509 22385 28543
rect 22385 28509 22419 28543
rect 22419 28509 22428 28543
rect 22376 28500 22428 28509
rect 23204 28500 23256 28552
rect 24308 28500 24360 28552
rect 23112 28364 23164 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3516 28203 3568 28212
rect 3516 28169 3525 28203
rect 3525 28169 3559 28203
rect 3559 28169 3568 28203
rect 3516 28160 3568 28169
rect 4620 28160 4672 28212
rect 5356 28160 5408 28212
rect 5540 28160 5592 28212
rect 7840 28203 7892 28212
rect 7840 28169 7865 28203
rect 7865 28169 7892 28203
rect 8024 28203 8076 28212
rect 7840 28160 7892 28169
rect 8024 28169 8033 28203
rect 8033 28169 8067 28203
rect 8067 28169 8076 28203
rect 8024 28160 8076 28169
rect 8668 28203 8720 28212
rect 8668 28169 8677 28203
rect 8677 28169 8711 28203
rect 8711 28169 8720 28203
rect 8668 28160 8720 28169
rect 9496 28203 9548 28212
rect 9496 28169 9505 28203
rect 9505 28169 9539 28203
rect 9539 28169 9548 28203
rect 9496 28160 9548 28169
rect 1676 28092 1728 28144
rect 6092 28092 6144 28144
rect 7656 28135 7708 28144
rect 7656 28101 7665 28135
rect 7665 28101 7699 28135
rect 7699 28101 7708 28135
rect 7656 28092 7708 28101
rect 2412 28067 2464 28076
rect 2412 28033 2446 28067
rect 2446 28033 2464 28067
rect 3976 28067 4028 28076
rect 2412 28024 2464 28033
rect 3976 28033 3985 28067
rect 3985 28033 4019 28067
rect 4019 28033 4028 28067
rect 3976 28024 4028 28033
rect 5632 28024 5684 28076
rect 5724 28067 5776 28076
rect 5724 28033 5733 28067
rect 5733 28033 5767 28067
rect 5767 28033 5776 28067
rect 9864 28092 9916 28144
rect 10508 28092 10560 28144
rect 5724 28024 5776 28033
rect 1584 27956 1636 28008
rect 2136 27999 2188 28008
rect 2136 27965 2145 27999
rect 2145 27965 2179 27999
rect 2179 27965 2188 27999
rect 2136 27956 2188 27965
rect 4804 27999 4856 28008
rect 4804 27965 4813 27999
rect 4813 27965 4847 27999
rect 4847 27965 4856 27999
rect 4804 27956 4856 27965
rect 5172 27999 5224 28008
rect 4712 27888 4764 27940
rect 5172 27965 5181 27999
rect 5181 27965 5215 27999
rect 5215 27965 5224 27999
rect 5172 27956 5224 27965
rect 8208 27956 8260 28008
rect 10416 28024 10468 28076
rect 10968 28024 11020 28076
rect 18696 28160 18748 28212
rect 18972 28203 19024 28212
rect 18972 28169 18981 28203
rect 18981 28169 19015 28203
rect 19015 28169 19024 28203
rect 18972 28160 19024 28169
rect 22192 28160 22244 28212
rect 14740 28092 14792 28144
rect 12900 28024 12952 28076
rect 14096 28024 14148 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 17132 28067 17184 28076
rect 17132 28033 17141 28067
rect 17141 28033 17175 28067
rect 17175 28033 17184 28067
rect 17132 28024 17184 28033
rect 18144 28024 18196 28076
rect 19340 28024 19392 28076
rect 20996 28092 21048 28144
rect 20536 28024 20588 28076
rect 21456 28024 21508 28076
rect 22100 28067 22152 28076
rect 22100 28033 22109 28067
rect 22109 28033 22143 28067
rect 22143 28033 22152 28067
rect 22100 28024 22152 28033
rect 22744 28024 22796 28076
rect 24216 28067 24268 28076
rect 24216 28033 24225 28067
rect 24225 28033 24259 28067
rect 24259 28033 24268 28067
rect 24216 28024 24268 28033
rect 24308 28067 24360 28076
rect 24308 28033 24317 28067
rect 24317 28033 24351 28067
rect 24351 28033 24360 28067
rect 24308 28024 24360 28033
rect 5264 27888 5316 27940
rect 5448 27820 5500 27872
rect 8484 27820 8536 27872
rect 9404 27956 9456 28008
rect 11796 27999 11848 28008
rect 11796 27965 11805 27999
rect 11805 27965 11839 27999
rect 11839 27965 11848 27999
rect 11796 27956 11848 27965
rect 12256 27999 12308 28008
rect 12256 27965 12265 27999
rect 12265 27965 12299 27999
rect 12299 27965 12308 27999
rect 12256 27956 12308 27965
rect 15568 27956 15620 28008
rect 16396 27956 16448 28008
rect 15476 27888 15528 27940
rect 18512 27888 18564 27940
rect 24400 27956 24452 28008
rect 24860 27956 24912 28008
rect 16212 27820 16264 27872
rect 16948 27820 17000 27872
rect 17408 27820 17460 27872
rect 18788 27863 18840 27872
rect 18788 27829 18797 27863
rect 18797 27829 18831 27863
rect 18831 27829 18840 27863
rect 18788 27820 18840 27829
rect 21180 27820 21232 27872
rect 21272 27820 21324 27872
rect 22652 27820 22704 27872
rect 24032 27863 24084 27872
rect 24032 27829 24041 27863
rect 24041 27829 24075 27863
rect 24075 27829 24084 27863
rect 24032 27820 24084 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2412 27616 2464 27668
rect 4804 27616 4856 27668
rect 4620 27548 4672 27600
rect 7840 27616 7892 27668
rect 10508 27616 10560 27668
rect 13636 27616 13688 27668
rect 16580 27616 16632 27668
rect 18512 27616 18564 27668
rect 18696 27616 18748 27668
rect 21272 27616 21324 27668
rect 5632 27548 5684 27600
rect 8300 27591 8352 27600
rect 8300 27557 8309 27591
rect 8309 27557 8343 27591
rect 8343 27557 8352 27591
rect 8300 27548 8352 27557
rect 12348 27548 12400 27600
rect 14556 27548 14608 27600
rect 1860 27412 1912 27464
rect 2688 27455 2740 27464
rect 2688 27421 2697 27455
rect 2697 27421 2731 27455
rect 2731 27421 2740 27455
rect 2688 27412 2740 27421
rect 4896 27480 4948 27532
rect 4620 27455 4672 27464
rect 4620 27421 4629 27455
rect 4629 27421 4663 27455
rect 4663 27421 4672 27455
rect 4620 27412 4672 27421
rect 5080 27412 5132 27464
rect 7840 27455 7892 27464
rect 3976 27344 4028 27396
rect 4988 27344 5040 27396
rect 7840 27421 7849 27455
rect 7849 27421 7883 27455
rect 7883 27421 7892 27455
rect 7840 27412 7892 27421
rect 5448 27344 5500 27396
rect 8208 27344 8260 27396
rect 11152 27480 11204 27532
rect 8576 27455 8628 27464
rect 8576 27421 8585 27455
rect 8585 27421 8619 27455
rect 8619 27421 8628 27455
rect 8576 27412 8628 27421
rect 11428 27412 11480 27464
rect 11980 27412 12032 27464
rect 9220 27344 9272 27396
rect 9312 27387 9364 27396
rect 9312 27353 9321 27387
rect 9321 27353 9355 27387
rect 9355 27353 9364 27387
rect 9312 27344 9364 27353
rect 9864 27344 9916 27396
rect 12256 27387 12308 27396
rect 12256 27353 12265 27387
rect 12265 27353 12299 27387
rect 12299 27353 12308 27387
rect 12256 27344 12308 27353
rect 12716 27480 12768 27532
rect 13084 27412 13136 27464
rect 13636 27480 13688 27532
rect 15016 27548 15068 27600
rect 15200 27548 15252 27600
rect 16212 27548 16264 27600
rect 18604 27548 18656 27600
rect 13728 27412 13780 27464
rect 14280 27412 14332 27464
rect 14832 27455 14884 27464
rect 14832 27421 14841 27455
rect 14841 27421 14875 27455
rect 14875 27421 14884 27455
rect 14832 27412 14884 27421
rect 13912 27344 13964 27396
rect 15016 27412 15068 27464
rect 15568 27480 15620 27532
rect 17040 27480 17092 27532
rect 17224 27523 17276 27532
rect 17224 27489 17233 27523
rect 17233 27489 17267 27523
rect 17267 27489 17276 27523
rect 17224 27480 17276 27489
rect 19432 27548 19484 27600
rect 20536 27548 20588 27600
rect 20720 27591 20772 27600
rect 20720 27557 20729 27591
rect 20729 27557 20763 27591
rect 20763 27557 20772 27591
rect 20720 27548 20772 27557
rect 25136 27591 25188 27600
rect 25136 27557 25145 27591
rect 25145 27557 25179 27591
rect 25179 27557 25188 27591
rect 25136 27548 25188 27557
rect 37832 27591 37884 27600
rect 37832 27557 37841 27591
rect 37841 27557 37875 27591
rect 37875 27557 37884 27591
rect 37832 27548 37884 27557
rect 20444 27523 20496 27532
rect 15476 27455 15528 27464
rect 15476 27421 15485 27455
rect 15485 27421 15519 27455
rect 15519 27421 15528 27455
rect 15476 27412 15528 27421
rect 16120 27412 16172 27464
rect 20444 27489 20453 27523
rect 20453 27489 20487 27523
rect 20487 27489 20496 27523
rect 20444 27480 20496 27489
rect 21548 27523 21600 27532
rect 21548 27489 21557 27523
rect 21557 27489 21591 27523
rect 21591 27489 21600 27523
rect 21548 27480 21600 27489
rect 17960 27455 18012 27464
rect 17960 27421 17969 27455
rect 17969 27421 18003 27455
rect 18003 27421 18012 27455
rect 17960 27412 18012 27421
rect 18144 27455 18196 27464
rect 18144 27421 18153 27455
rect 18153 27421 18187 27455
rect 18187 27421 18196 27455
rect 18144 27412 18196 27421
rect 18236 27455 18288 27464
rect 18236 27421 18245 27455
rect 18245 27421 18279 27455
rect 18279 27421 18288 27455
rect 18236 27412 18288 27421
rect 1768 27319 1820 27328
rect 1768 27285 1777 27319
rect 1777 27285 1811 27319
rect 1811 27285 1820 27319
rect 1768 27276 1820 27285
rect 8392 27276 8444 27328
rect 10508 27319 10560 27328
rect 10508 27285 10517 27319
rect 10517 27285 10551 27319
rect 10551 27285 10560 27319
rect 10508 27276 10560 27285
rect 11336 27319 11388 27328
rect 11336 27285 11345 27319
rect 11345 27285 11379 27319
rect 11379 27285 11388 27319
rect 11336 27276 11388 27285
rect 12072 27276 12124 27328
rect 12440 27319 12492 27328
rect 12440 27285 12449 27319
rect 12449 27285 12483 27319
rect 12483 27285 12492 27319
rect 12440 27276 12492 27285
rect 14280 27276 14332 27328
rect 14556 27276 14608 27328
rect 16948 27344 17000 27396
rect 15384 27276 15436 27328
rect 17592 27344 17644 27396
rect 17132 27276 17184 27328
rect 18236 27276 18288 27328
rect 18420 27319 18472 27328
rect 18420 27285 18429 27319
rect 18429 27285 18463 27319
rect 18463 27285 18472 27319
rect 18420 27276 18472 27285
rect 19340 27344 19392 27396
rect 23480 27480 23532 27532
rect 25044 27480 25096 27532
rect 22652 27412 22704 27464
rect 24032 27412 24084 27464
rect 38016 27455 38068 27464
rect 38016 27421 38025 27455
rect 38025 27421 38059 27455
rect 38059 27421 38068 27455
rect 38016 27412 38068 27421
rect 24860 27344 24912 27396
rect 20996 27276 21048 27328
rect 22100 27276 22152 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 1860 27115 1912 27124
rect 1860 27081 1869 27115
rect 1869 27081 1903 27115
rect 1903 27081 1912 27115
rect 1860 27072 1912 27081
rect 5356 27072 5408 27124
rect 7840 27072 7892 27124
rect 9312 27072 9364 27124
rect 11980 27115 12032 27124
rect 11980 27081 11989 27115
rect 11989 27081 12023 27115
rect 12023 27081 12032 27115
rect 11980 27072 12032 27081
rect 12072 27072 12124 27124
rect 14280 27115 14332 27124
rect 14280 27081 14289 27115
rect 14289 27081 14323 27115
rect 14323 27081 14332 27115
rect 14280 27072 14332 27081
rect 2044 26979 2096 26988
rect 2044 26945 2053 26979
rect 2053 26945 2087 26979
rect 2087 26945 2096 26979
rect 2044 26936 2096 26945
rect 3516 26979 3568 26988
rect 3516 26945 3525 26979
rect 3525 26945 3559 26979
rect 3559 26945 3568 26979
rect 3516 26936 3568 26945
rect 3608 26979 3660 26988
rect 3608 26945 3617 26979
rect 3617 26945 3651 26979
rect 3651 26945 3660 26979
rect 4712 27004 4764 27056
rect 3608 26936 3660 26945
rect 4988 26936 5040 26988
rect 5172 27004 5224 27056
rect 5540 27004 5592 27056
rect 5264 26979 5316 26988
rect 5264 26945 5273 26979
rect 5273 26945 5307 26979
rect 5307 26945 5316 26979
rect 5264 26936 5316 26945
rect 5356 26979 5408 26988
rect 5356 26945 5365 26979
rect 5365 26945 5399 26979
rect 5399 26945 5408 26979
rect 5816 26979 5868 26988
rect 5356 26936 5408 26945
rect 5816 26945 5825 26979
rect 5825 26945 5859 26979
rect 5859 26945 5868 26979
rect 5816 26936 5868 26945
rect 6460 27004 6512 27056
rect 11336 27004 11388 27056
rect 12716 27004 12768 27056
rect 13912 27004 13964 27056
rect 6184 26936 6236 26988
rect 8208 26936 8260 26988
rect 9404 26936 9456 26988
rect 13636 26979 13688 26988
rect 3884 26868 3936 26920
rect 3332 26775 3384 26784
rect 3332 26741 3341 26775
rect 3341 26741 3375 26775
rect 3375 26741 3384 26775
rect 3332 26732 3384 26741
rect 4804 26800 4856 26852
rect 7748 26800 7800 26852
rect 8668 26911 8720 26920
rect 8668 26877 8677 26911
rect 8677 26877 8711 26911
rect 8711 26877 8720 26911
rect 8668 26868 8720 26877
rect 9588 26868 9640 26920
rect 9680 26868 9732 26920
rect 4620 26732 4672 26784
rect 4896 26775 4948 26784
rect 4896 26741 4905 26775
rect 4905 26741 4939 26775
rect 4939 26741 4948 26775
rect 4896 26732 4948 26741
rect 5908 26775 5960 26784
rect 5908 26741 5917 26775
rect 5917 26741 5951 26775
rect 5951 26741 5960 26775
rect 5908 26732 5960 26741
rect 13636 26945 13645 26979
rect 13645 26945 13679 26979
rect 13679 26945 13688 26979
rect 13636 26936 13688 26945
rect 13728 26936 13780 26988
rect 14464 27004 14516 27056
rect 15568 27072 15620 27124
rect 17408 27072 17460 27124
rect 17960 27072 18012 27124
rect 15200 26936 15252 26988
rect 15476 26936 15528 26988
rect 18420 27004 18472 27056
rect 19340 27072 19392 27124
rect 24216 27072 24268 27124
rect 16488 26936 16540 26988
rect 16948 26979 17000 26988
rect 15660 26868 15712 26920
rect 16120 26868 16172 26920
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 18236 26936 18288 26988
rect 18972 26936 19024 26988
rect 24952 27004 25004 27056
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 23848 26979 23900 26988
rect 13268 26732 13320 26784
rect 16396 26800 16448 26852
rect 14832 26732 14884 26784
rect 15476 26732 15528 26784
rect 15936 26775 15988 26784
rect 15936 26741 15945 26775
rect 15945 26741 15979 26775
rect 15979 26741 15988 26775
rect 15936 26732 15988 26741
rect 16120 26775 16172 26784
rect 16120 26741 16129 26775
rect 16129 26741 16163 26775
rect 16163 26741 16172 26775
rect 16856 26800 16908 26852
rect 17684 26800 17736 26852
rect 18144 26868 18196 26920
rect 18880 26911 18932 26920
rect 18420 26800 18472 26852
rect 16120 26732 16172 26741
rect 17500 26732 17552 26784
rect 18880 26877 18889 26911
rect 18889 26877 18923 26911
rect 18923 26877 18932 26911
rect 18880 26868 18932 26877
rect 23848 26945 23857 26979
rect 23857 26945 23891 26979
rect 23891 26945 23900 26979
rect 23848 26936 23900 26945
rect 23112 26868 23164 26920
rect 24400 26979 24452 26988
rect 24400 26945 24409 26979
rect 24409 26945 24443 26979
rect 24443 26945 24452 26979
rect 24400 26936 24452 26945
rect 24860 26936 24912 26988
rect 19892 26800 19944 26852
rect 22284 26800 22336 26852
rect 38016 26800 38068 26852
rect 22192 26732 22244 26784
rect 24768 26732 24820 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3976 26571 4028 26580
rect 3976 26537 3985 26571
rect 3985 26537 4019 26571
rect 4019 26537 4028 26571
rect 3976 26528 4028 26537
rect 5448 26528 5500 26580
rect 6184 26571 6236 26580
rect 6184 26537 6193 26571
rect 6193 26537 6227 26571
rect 6227 26537 6236 26571
rect 6184 26528 6236 26537
rect 9220 26528 9272 26580
rect 12256 26571 12308 26580
rect 3516 26460 3568 26512
rect 5080 26460 5132 26512
rect 5540 26460 5592 26512
rect 5172 26392 5224 26444
rect 5908 26392 5960 26444
rect 7748 26435 7800 26444
rect 1584 26324 1636 26376
rect 3884 26324 3936 26376
rect 4160 26367 4212 26376
rect 4160 26333 4166 26367
rect 4166 26333 4200 26367
rect 4200 26333 4212 26367
rect 4160 26324 4212 26333
rect 4620 26367 4672 26376
rect 4620 26333 4629 26367
rect 4629 26333 4663 26367
rect 4663 26333 4672 26367
rect 5080 26367 5132 26376
rect 4620 26324 4672 26333
rect 5080 26333 5089 26367
rect 5089 26333 5123 26367
rect 5123 26333 5132 26367
rect 5080 26324 5132 26333
rect 6460 26367 6512 26376
rect 6460 26333 6469 26367
rect 6469 26333 6503 26367
rect 6503 26333 6512 26367
rect 6460 26324 6512 26333
rect 7748 26401 7757 26435
rect 7757 26401 7791 26435
rect 7791 26401 7800 26435
rect 7748 26392 7800 26401
rect 8576 26392 8628 26444
rect 12256 26537 12265 26571
rect 12265 26537 12299 26571
rect 12299 26537 12308 26571
rect 12256 26528 12308 26537
rect 13084 26571 13136 26580
rect 13084 26537 13093 26571
rect 13093 26537 13127 26571
rect 13127 26537 13136 26571
rect 13084 26528 13136 26537
rect 14556 26528 14608 26580
rect 14924 26571 14976 26580
rect 14924 26537 14933 26571
rect 14933 26537 14967 26571
rect 14967 26537 14976 26571
rect 14924 26528 14976 26537
rect 15568 26528 15620 26580
rect 15844 26528 15896 26580
rect 18052 26571 18104 26580
rect 18052 26537 18061 26571
rect 18061 26537 18095 26571
rect 18095 26537 18104 26571
rect 18328 26571 18380 26580
rect 18052 26528 18104 26537
rect 18328 26537 18337 26571
rect 18337 26537 18371 26571
rect 18371 26537 18380 26571
rect 18328 26528 18380 26537
rect 18880 26528 18932 26580
rect 25044 26571 25096 26580
rect 6828 26367 6880 26376
rect 2596 26256 2648 26308
rect 3608 26256 3660 26308
rect 4436 26256 4488 26308
rect 5724 26256 5776 26308
rect 6828 26333 6837 26367
rect 6837 26333 6871 26367
rect 6871 26333 6880 26367
rect 6828 26324 6880 26333
rect 7288 26256 7340 26308
rect 8392 26256 8444 26308
rect 9588 26324 9640 26376
rect 5356 26188 5408 26240
rect 8024 26188 8076 26240
rect 9772 26299 9824 26308
rect 9772 26265 9806 26299
rect 9806 26265 9824 26299
rect 14464 26392 14516 26444
rect 13728 26367 13780 26376
rect 13728 26333 13737 26367
rect 13737 26333 13771 26367
rect 13771 26333 13780 26367
rect 13728 26324 13780 26333
rect 17040 26503 17092 26512
rect 16120 26392 16172 26444
rect 15384 26367 15436 26376
rect 15384 26333 15393 26367
rect 15393 26333 15427 26367
rect 15427 26333 15436 26367
rect 15384 26324 15436 26333
rect 9772 26256 9824 26265
rect 12072 26256 12124 26308
rect 12900 26299 12952 26308
rect 12900 26265 12909 26299
rect 12909 26265 12943 26299
rect 12943 26265 12952 26299
rect 12900 26256 12952 26265
rect 13452 26256 13504 26308
rect 9680 26188 9732 26240
rect 14556 26256 14608 26308
rect 15936 26324 15988 26376
rect 17040 26469 17049 26503
rect 17049 26469 17083 26503
rect 17083 26469 17092 26503
rect 17040 26460 17092 26469
rect 20536 26460 20588 26512
rect 22100 26460 22152 26512
rect 23480 26503 23532 26512
rect 23480 26469 23489 26503
rect 23489 26469 23523 26503
rect 23523 26469 23532 26503
rect 23480 26460 23532 26469
rect 19340 26392 19392 26444
rect 16028 26299 16080 26308
rect 16028 26265 16037 26299
rect 16037 26265 16071 26299
rect 16071 26265 16080 26299
rect 16028 26256 16080 26265
rect 17316 26256 17368 26308
rect 18236 26324 18288 26376
rect 18420 26324 18472 26376
rect 20076 26392 20128 26444
rect 20352 26392 20404 26444
rect 19892 26324 19944 26376
rect 20996 26367 21048 26376
rect 20996 26333 21005 26367
rect 21005 26333 21039 26367
rect 21039 26333 21048 26367
rect 20996 26324 21048 26333
rect 25044 26537 25053 26571
rect 25053 26537 25087 26571
rect 25087 26537 25096 26571
rect 25044 26528 25096 26537
rect 19248 26188 19300 26240
rect 22192 26256 22244 26308
rect 24768 26367 24820 26376
rect 24768 26333 24777 26367
rect 24777 26333 24811 26367
rect 24811 26333 24820 26367
rect 24768 26324 24820 26333
rect 37188 26324 37240 26376
rect 37740 26367 37792 26376
rect 37740 26333 37749 26367
rect 37749 26333 37783 26367
rect 37783 26333 37792 26367
rect 37740 26324 37792 26333
rect 21732 26188 21784 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2596 26027 2648 26036
rect 2596 25993 2605 26027
rect 2605 25993 2639 26027
rect 2639 25993 2648 26027
rect 2596 25984 2648 25993
rect 4620 25984 4672 26036
rect 4804 25984 4856 26036
rect 3332 25916 3384 25968
rect 4528 25916 4580 25968
rect 2688 25891 2740 25900
rect 2688 25857 2697 25891
rect 2697 25857 2731 25891
rect 2731 25857 2740 25891
rect 2688 25848 2740 25857
rect 4068 25891 4120 25900
rect 4068 25857 4077 25891
rect 4077 25857 4111 25891
rect 4111 25857 4120 25891
rect 4068 25848 4120 25857
rect 4988 25712 5040 25764
rect 5264 25916 5316 25968
rect 5540 25891 5592 25900
rect 5540 25857 5549 25891
rect 5549 25857 5583 25891
rect 5583 25857 5592 25891
rect 5540 25848 5592 25857
rect 9864 25984 9916 26036
rect 12440 25984 12492 26036
rect 5356 25780 5408 25832
rect 6460 25848 6512 25900
rect 6736 25891 6788 25900
rect 6736 25857 6745 25891
rect 6745 25857 6779 25891
rect 6779 25857 6788 25891
rect 6736 25848 6788 25857
rect 6644 25780 6696 25832
rect 7104 25848 7156 25900
rect 7472 25891 7524 25900
rect 7472 25857 7481 25891
rect 7481 25857 7515 25891
rect 7515 25857 7524 25891
rect 7472 25848 7524 25857
rect 7656 25891 7708 25900
rect 7656 25857 7665 25891
rect 7665 25857 7699 25891
rect 7699 25857 7708 25891
rect 7656 25848 7708 25857
rect 8576 25848 8628 25900
rect 10508 25916 10560 25968
rect 8852 25848 8904 25900
rect 9680 25891 9732 25900
rect 9680 25857 9689 25891
rect 9689 25857 9723 25891
rect 9723 25857 9732 25891
rect 9680 25848 9732 25857
rect 12072 25891 12124 25900
rect 8760 25823 8812 25832
rect 8760 25789 8769 25823
rect 8769 25789 8803 25823
rect 8803 25789 8812 25823
rect 8760 25780 8812 25789
rect 12072 25857 12081 25891
rect 12081 25857 12115 25891
rect 12115 25857 12124 25891
rect 12072 25848 12124 25857
rect 12900 25848 12952 25900
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 13636 25848 13688 25900
rect 15200 25984 15252 26036
rect 18972 26027 19024 26036
rect 18972 25993 18981 26027
rect 18981 25993 19015 26027
rect 19015 25993 19024 26027
rect 18972 25984 19024 25993
rect 20444 25984 20496 26036
rect 23848 25984 23900 26036
rect 24952 26027 25004 26036
rect 24952 25993 24961 26027
rect 24961 25993 24995 26027
rect 24995 25993 25004 26027
rect 24952 25984 25004 25993
rect 16028 25916 16080 25968
rect 18144 25916 18196 25968
rect 18604 25916 18656 25968
rect 19248 25959 19300 25968
rect 19248 25925 19257 25959
rect 19257 25925 19291 25959
rect 19291 25925 19300 25959
rect 19248 25916 19300 25925
rect 20168 25916 20220 25968
rect 14832 25891 14884 25900
rect 14832 25857 14841 25891
rect 14841 25857 14875 25891
rect 14875 25857 14884 25891
rect 14832 25848 14884 25857
rect 15016 25891 15068 25900
rect 15016 25857 15025 25891
rect 15025 25857 15059 25891
rect 15059 25857 15068 25891
rect 15016 25848 15068 25857
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 17316 25848 17368 25900
rect 19156 25891 19208 25900
rect 19156 25857 19165 25891
rect 19165 25857 19199 25891
rect 19199 25857 19208 25891
rect 19156 25848 19208 25857
rect 19892 25848 19944 25900
rect 20076 25891 20128 25900
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 20260 25891 20312 25900
rect 20260 25857 20269 25891
rect 20269 25857 20303 25891
rect 20303 25857 20312 25891
rect 20260 25848 20312 25857
rect 20996 25891 21048 25900
rect 20996 25857 21005 25891
rect 21005 25857 21039 25891
rect 21039 25857 21048 25891
rect 22468 25891 22520 25900
rect 20996 25848 21048 25857
rect 5724 25712 5776 25764
rect 19524 25780 19576 25832
rect 19708 25780 19760 25832
rect 19984 25780 20036 25832
rect 20628 25780 20680 25832
rect 22468 25857 22477 25891
rect 22477 25857 22511 25891
rect 22511 25857 22520 25891
rect 22468 25848 22520 25857
rect 23480 25848 23532 25900
rect 24400 25848 24452 25900
rect 22744 25780 22796 25832
rect 23296 25780 23348 25832
rect 9772 25712 9824 25764
rect 9864 25712 9916 25764
rect 24676 25780 24728 25832
rect 4896 25687 4948 25696
rect 4896 25653 4905 25687
rect 4905 25653 4939 25687
rect 4939 25653 4948 25687
rect 4896 25644 4948 25653
rect 7012 25644 7064 25696
rect 7564 25644 7616 25696
rect 8300 25644 8352 25696
rect 10048 25644 10100 25696
rect 13176 25644 13228 25696
rect 13636 25687 13688 25696
rect 13636 25653 13645 25687
rect 13645 25653 13679 25687
rect 13679 25653 13688 25687
rect 13636 25644 13688 25653
rect 14372 25644 14424 25696
rect 14648 25644 14700 25696
rect 15292 25644 15344 25696
rect 16856 25644 16908 25696
rect 17684 25644 17736 25696
rect 20076 25687 20128 25696
rect 20076 25653 20085 25687
rect 20085 25653 20119 25687
rect 20119 25653 20128 25687
rect 20076 25644 20128 25653
rect 22652 25687 22704 25696
rect 22652 25653 22661 25687
rect 22661 25653 22695 25687
rect 22695 25653 22704 25687
rect 22652 25644 22704 25653
rect 23756 25687 23808 25696
rect 23756 25653 23765 25687
rect 23765 25653 23799 25687
rect 23799 25653 23808 25687
rect 23756 25644 23808 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4068 25440 4120 25492
rect 6736 25440 6788 25492
rect 8392 25483 8444 25492
rect 8392 25449 8401 25483
rect 8401 25449 8435 25483
rect 8435 25449 8444 25483
rect 8392 25440 8444 25449
rect 8576 25483 8628 25492
rect 8576 25449 8585 25483
rect 8585 25449 8619 25483
rect 8619 25449 8628 25483
rect 8576 25440 8628 25449
rect 9680 25440 9732 25492
rect 13360 25440 13412 25492
rect 15844 25440 15896 25492
rect 19156 25440 19208 25492
rect 5632 25372 5684 25424
rect 4712 25236 4764 25288
rect 4804 25279 4856 25288
rect 4804 25245 4813 25279
rect 4813 25245 4847 25279
rect 4847 25245 4856 25279
rect 4804 25236 4856 25245
rect 5908 25372 5960 25424
rect 6092 25372 6144 25424
rect 9864 25372 9916 25424
rect 17868 25372 17920 25424
rect 6828 25236 6880 25288
rect 7196 25236 7248 25288
rect 7564 25279 7616 25288
rect 7564 25245 7573 25279
rect 7573 25245 7607 25279
rect 7607 25245 7616 25279
rect 7564 25236 7616 25245
rect 5356 25168 5408 25220
rect 5264 25143 5316 25152
rect 5264 25109 5273 25143
rect 5273 25109 5307 25143
rect 5307 25109 5316 25143
rect 5264 25100 5316 25109
rect 6460 25211 6512 25220
rect 6460 25177 6469 25211
rect 6469 25177 6503 25211
rect 6503 25177 6512 25211
rect 6460 25168 6512 25177
rect 8668 25236 8720 25288
rect 8484 25168 8536 25220
rect 9220 25236 9272 25288
rect 9956 25279 10008 25288
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 9956 25236 10008 25245
rect 10508 25236 10560 25288
rect 6092 25100 6144 25152
rect 6644 25143 6696 25152
rect 6644 25109 6669 25143
rect 6669 25109 6696 25143
rect 6644 25100 6696 25109
rect 7104 25100 7156 25152
rect 7288 25100 7340 25152
rect 10692 25168 10744 25220
rect 11888 25168 11940 25220
rect 12716 25168 12768 25220
rect 16120 25304 16172 25356
rect 16488 25304 16540 25356
rect 17408 25347 17460 25356
rect 17408 25313 17417 25347
rect 17417 25313 17451 25347
rect 17451 25313 17460 25347
rect 17408 25304 17460 25313
rect 14556 25236 14608 25288
rect 14372 25168 14424 25220
rect 16028 25236 16080 25288
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 18512 25304 18564 25356
rect 18880 25372 18932 25424
rect 19340 25372 19392 25424
rect 20536 25440 20588 25492
rect 23020 25440 23072 25492
rect 21732 25415 21784 25424
rect 21732 25381 21741 25415
rect 21741 25381 21775 25415
rect 21775 25381 21784 25415
rect 21732 25372 21784 25381
rect 22468 25372 22520 25424
rect 18880 25279 18932 25288
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 18880 25236 18932 25245
rect 19984 25236 20036 25288
rect 22836 25347 22888 25356
rect 22836 25313 22845 25347
rect 22845 25313 22879 25347
rect 22879 25313 22888 25347
rect 22836 25304 22888 25313
rect 19340 25168 19392 25220
rect 19708 25168 19760 25220
rect 10140 25143 10192 25152
rect 10140 25109 10149 25143
rect 10149 25109 10183 25143
rect 10183 25109 10192 25143
rect 10140 25100 10192 25109
rect 10968 25143 11020 25152
rect 10968 25109 10977 25143
rect 10977 25109 11011 25143
rect 11011 25109 11020 25143
rect 10968 25100 11020 25109
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 14924 25143 14976 25152
rect 14924 25109 14933 25143
rect 14933 25109 14967 25143
rect 14967 25109 14976 25143
rect 14924 25100 14976 25109
rect 15384 25100 15436 25152
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 17316 25100 17368 25152
rect 17960 25100 18012 25152
rect 18696 25100 18748 25152
rect 18880 25100 18932 25152
rect 20720 25100 20772 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 5264 24828 5316 24880
rect 2320 24760 2372 24812
rect 2412 24803 2464 24812
rect 2412 24769 2421 24803
rect 2421 24769 2455 24803
rect 2455 24769 2464 24803
rect 2412 24760 2464 24769
rect 2688 24760 2740 24812
rect 3148 24803 3200 24812
rect 3148 24769 3157 24803
rect 3157 24769 3191 24803
rect 3191 24769 3200 24803
rect 3148 24760 3200 24769
rect 6460 24760 6512 24812
rect 7932 24760 7984 24812
rect 10140 24828 10192 24880
rect 10968 24828 11020 24880
rect 14372 24871 14424 24880
rect 14372 24837 14381 24871
rect 14381 24837 14415 24871
rect 14415 24837 14424 24871
rect 14372 24828 14424 24837
rect 15752 24896 15804 24948
rect 18880 24896 18932 24948
rect 19340 24939 19392 24948
rect 19340 24905 19349 24939
rect 19349 24905 19383 24939
rect 19383 24905 19392 24939
rect 19340 24896 19392 24905
rect 9956 24760 10008 24812
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 1584 24692 1636 24744
rect 8024 24735 8076 24744
rect 8024 24701 8033 24735
rect 8033 24701 8067 24735
rect 8067 24701 8076 24735
rect 8024 24692 8076 24701
rect 6000 24667 6052 24676
rect 6000 24633 6009 24667
rect 6009 24633 6043 24667
rect 6043 24633 6052 24667
rect 6000 24624 6052 24633
rect 2228 24599 2280 24608
rect 2228 24565 2237 24599
rect 2237 24565 2271 24599
rect 2271 24565 2280 24599
rect 2228 24556 2280 24565
rect 3056 24556 3108 24608
rect 3608 24599 3660 24608
rect 3608 24565 3617 24599
rect 3617 24565 3651 24599
rect 3651 24565 3660 24599
rect 3608 24556 3660 24565
rect 4896 24556 4948 24608
rect 5264 24556 5316 24608
rect 10048 24692 10100 24744
rect 10692 24760 10744 24812
rect 11888 24803 11940 24812
rect 11888 24769 11897 24803
rect 11897 24769 11931 24803
rect 11931 24769 11940 24803
rect 11888 24760 11940 24769
rect 12716 24760 12768 24812
rect 14556 24803 14608 24812
rect 14556 24769 14565 24803
rect 14565 24769 14599 24803
rect 14599 24769 14608 24803
rect 14556 24760 14608 24769
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 9772 24624 9824 24676
rect 10692 24624 10744 24676
rect 13360 24692 13412 24744
rect 13636 24692 13688 24744
rect 9680 24556 9732 24608
rect 10600 24556 10652 24608
rect 11796 24556 11848 24608
rect 16120 24760 16172 24812
rect 17500 24803 17552 24812
rect 17500 24769 17509 24803
rect 17509 24769 17543 24803
rect 17543 24769 17552 24803
rect 17500 24760 17552 24769
rect 17960 24828 18012 24880
rect 17684 24806 17736 24812
rect 17684 24772 17693 24806
rect 17693 24772 17727 24806
rect 17727 24772 17736 24806
rect 17684 24760 17736 24772
rect 17868 24803 17920 24812
rect 17868 24769 17877 24803
rect 17877 24769 17911 24803
rect 17911 24769 17920 24803
rect 17868 24760 17920 24769
rect 18880 24760 18932 24812
rect 19248 24760 19300 24812
rect 20260 24896 20312 24948
rect 20720 24896 20772 24948
rect 18788 24624 18840 24676
rect 19340 24692 19392 24744
rect 20076 24828 20128 24880
rect 19800 24692 19852 24744
rect 19708 24624 19760 24676
rect 20536 24760 20588 24812
rect 22652 24828 22704 24880
rect 22836 24896 22888 24948
rect 23388 24896 23440 24948
rect 24768 24871 24820 24880
rect 24768 24837 24777 24871
rect 24777 24837 24811 24871
rect 24811 24837 24820 24871
rect 24768 24828 24820 24837
rect 22054 24760 22106 24812
rect 24584 24803 24636 24812
rect 20168 24624 20220 24676
rect 22100 24624 22152 24676
rect 24584 24769 24593 24803
rect 24593 24769 24627 24803
rect 24627 24769 24636 24803
rect 24584 24760 24636 24769
rect 19156 24556 19208 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2320 24352 2372 24404
rect 7012 24352 7064 24404
rect 7932 24395 7984 24404
rect 7932 24361 7941 24395
rect 7941 24361 7975 24395
rect 7975 24361 7984 24395
rect 7932 24352 7984 24361
rect 10232 24352 10284 24404
rect 14188 24352 14240 24404
rect 19708 24395 19760 24404
rect 3424 24284 3476 24336
rect 1584 24259 1636 24268
rect 1584 24225 1593 24259
rect 1593 24225 1627 24259
rect 1627 24225 1636 24259
rect 1584 24216 1636 24225
rect 4896 24216 4948 24268
rect 6000 24259 6052 24268
rect 6000 24225 6009 24259
rect 6009 24225 6043 24259
rect 6043 24225 6052 24259
rect 6000 24216 6052 24225
rect 7012 24216 7064 24268
rect 8760 24284 8812 24336
rect 19708 24361 19717 24395
rect 19717 24361 19751 24395
rect 19751 24361 19760 24395
rect 19708 24352 19760 24361
rect 20444 24352 20496 24404
rect 20904 24395 20956 24404
rect 20904 24361 20913 24395
rect 20913 24361 20947 24395
rect 20947 24361 20956 24395
rect 20904 24352 20956 24361
rect 20076 24284 20128 24336
rect 8024 24216 8076 24268
rect 2228 24148 2280 24200
rect 3148 24148 3200 24200
rect 4436 24148 4488 24200
rect 4620 24191 4672 24200
rect 4620 24157 4629 24191
rect 4629 24157 4663 24191
rect 4663 24157 4672 24191
rect 6092 24191 6144 24200
rect 4620 24148 4672 24157
rect 6092 24157 6101 24191
rect 6101 24157 6135 24191
rect 6135 24157 6144 24191
rect 6092 24148 6144 24157
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 6000 24080 6052 24132
rect 6736 24080 6788 24132
rect 4528 24012 4580 24064
rect 5356 24012 5408 24064
rect 7288 24012 7340 24064
rect 9956 24148 10008 24200
rect 13452 24191 13504 24200
rect 8852 24080 8904 24132
rect 10508 24080 10560 24132
rect 13452 24157 13461 24191
rect 13461 24157 13495 24191
rect 13495 24157 13504 24191
rect 13452 24148 13504 24157
rect 12164 24080 12216 24132
rect 12992 24080 13044 24132
rect 8116 24055 8168 24064
rect 8116 24021 8125 24055
rect 8125 24021 8159 24055
rect 8159 24021 8168 24055
rect 8116 24012 8168 24021
rect 8208 24012 8260 24064
rect 13268 24055 13320 24064
rect 13268 24021 13277 24055
rect 13277 24021 13311 24055
rect 13311 24021 13320 24055
rect 13268 24012 13320 24021
rect 14096 24148 14148 24200
rect 19156 24216 19208 24268
rect 14924 24080 14976 24132
rect 16396 24191 16448 24200
rect 16396 24157 16405 24191
rect 16405 24157 16439 24191
rect 16439 24157 16448 24191
rect 16396 24148 16448 24157
rect 16580 24191 16632 24200
rect 16580 24157 16589 24191
rect 16589 24157 16623 24191
rect 16623 24157 16632 24191
rect 16580 24148 16632 24157
rect 17500 24148 17552 24200
rect 20352 24148 20404 24200
rect 20536 24191 20588 24200
rect 20536 24157 20545 24191
rect 20545 24157 20579 24191
rect 20579 24157 20588 24191
rect 20536 24148 20588 24157
rect 22100 24352 22152 24404
rect 22376 24352 22428 24404
rect 23756 24216 23808 24268
rect 23388 24148 23440 24200
rect 19340 24080 19392 24132
rect 21272 24080 21324 24132
rect 23480 24080 23532 24132
rect 15660 24055 15712 24064
rect 15660 24021 15669 24055
rect 15669 24021 15703 24055
rect 15703 24021 15712 24055
rect 15660 24012 15712 24021
rect 16304 24012 16356 24064
rect 16764 24012 16816 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3240 23808 3292 23860
rect 3700 23808 3752 23860
rect 6000 23851 6052 23860
rect 6000 23817 6009 23851
rect 6009 23817 6043 23851
rect 6043 23817 6052 23851
rect 6000 23808 6052 23817
rect 6092 23808 6144 23860
rect 8116 23808 8168 23860
rect 9772 23851 9824 23860
rect 9772 23817 9781 23851
rect 9781 23817 9815 23851
rect 9815 23817 9824 23851
rect 9772 23808 9824 23817
rect 12164 23851 12216 23860
rect 12164 23817 12173 23851
rect 12173 23817 12207 23851
rect 12207 23817 12216 23851
rect 12164 23808 12216 23817
rect 3608 23740 3660 23792
rect 3240 23672 3292 23724
rect 4712 23672 4764 23724
rect 8208 23740 8260 23792
rect 3424 23647 3476 23656
rect 3424 23613 3433 23647
rect 3433 23613 3467 23647
rect 3467 23613 3476 23647
rect 3424 23604 3476 23613
rect 4620 23604 4672 23656
rect 7288 23672 7340 23724
rect 9680 23740 9732 23792
rect 14188 23808 14240 23860
rect 14280 23851 14332 23860
rect 14280 23817 14289 23851
rect 14289 23817 14323 23851
rect 14323 23817 14332 23851
rect 14280 23808 14332 23817
rect 14924 23851 14976 23860
rect 8668 23715 8720 23724
rect 8668 23681 8702 23715
rect 8702 23681 8720 23715
rect 8668 23672 8720 23681
rect 12532 23672 12584 23724
rect 8024 23604 8076 23656
rect 12808 23672 12860 23724
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 13360 23715 13412 23724
rect 13360 23681 13369 23715
rect 13369 23681 13403 23715
rect 13403 23681 13412 23715
rect 13360 23672 13412 23681
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 16212 23851 16264 23860
rect 16212 23817 16221 23851
rect 16221 23817 16255 23851
rect 16255 23817 16264 23851
rect 16212 23808 16264 23817
rect 16488 23808 16540 23860
rect 18236 23851 18288 23860
rect 18236 23817 18245 23851
rect 18245 23817 18279 23851
rect 18279 23817 18288 23851
rect 18236 23808 18288 23817
rect 20720 23808 20772 23860
rect 23388 23808 23440 23860
rect 16028 23715 16080 23724
rect 16028 23681 16037 23715
rect 16037 23681 16071 23715
rect 16071 23681 16080 23715
rect 16028 23672 16080 23681
rect 16304 23715 16356 23724
rect 16304 23681 16313 23715
rect 16313 23681 16347 23715
rect 16347 23681 16356 23715
rect 16304 23672 16356 23681
rect 4436 23511 4488 23520
rect 4436 23477 4445 23511
rect 4445 23477 4479 23511
rect 4479 23477 4488 23511
rect 4436 23468 4488 23477
rect 4804 23468 4856 23520
rect 13452 23604 13504 23656
rect 20996 23740 21048 23792
rect 22008 23783 22060 23792
rect 22008 23749 22017 23783
rect 22017 23749 22051 23783
rect 22051 23749 22060 23783
rect 22008 23740 22060 23749
rect 11888 23536 11940 23588
rect 13912 23579 13964 23588
rect 13912 23545 13921 23579
rect 13921 23545 13955 23579
rect 13955 23545 13964 23579
rect 13912 23536 13964 23545
rect 14096 23536 14148 23588
rect 11152 23511 11204 23520
rect 11152 23477 11161 23511
rect 11161 23477 11195 23511
rect 11195 23477 11204 23511
rect 11152 23468 11204 23477
rect 13268 23468 13320 23520
rect 20536 23672 20588 23724
rect 23204 23715 23256 23724
rect 18696 23647 18748 23656
rect 18696 23613 18705 23647
rect 18705 23613 18739 23647
rect 18739 23613 18748 23647
rect 18696 23604 18748 23613
rect 19156 23604 19208 23656
rect 19340 23604 19392 23656
rect 21272 23604 21324 23656
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 23296 23672 23348 23724
rect 23940 23672 23992 23724
rect 22468 23536 22520 23588
rect 23480 23536 23532 23588
rect 20996 23468 21048 23520
rect 22376 23511 22428 23520
rect 22376 23477 22385 23511
rect 22385 23477 22419 23511
rect 22419 23477 22428 23511
rect 22376 23468 22428 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8668 23264 8720 23316
rect 8852 23264 8904 23316
rect 12808 23264 12860 23316
rect 16028 23264 16080 23316
rect 18144 23264 18196 23316
rect 18604 23264 18656 23316
rect 19432 23264 19484 23316
rect 20904 23307 20956 23316
rect 20904 23273 20913 23307
rect 20913 23273 20947 23307
rect 20947 23273 20956 23307
rect 20904 23264 20956 23273
rect 23940 23307 23992 23316
rect 23940 23273 23949 23307
rect 23949 23273 23983 23307
rect 23983 23273 23992 23307
rect 23940 23264 23992 23273
rect 4804 23196 4856 23248
rect 6552 23239 6604 23248
rect 6552 23205 6561 23239
rect 6561 23205 6595 23239
rect 6595 23205 6604 23239
rect 6552 23196 6604 23205
rect 4344 23128 4396 23180
rect 4712 23128 4764 23180
rect 5172 23128 5224 23180
rect 15384 23171 15436 23180
rect 5356 23060 5408 23112
rect 6092 23103 6144 23112
rect 6092 23069 6101 23103
rect 6101 23069 6135 23103
rect 6135 23069 6144 23103
rect 6092 23060 6144 23069
rect 7104 23060 7156 23112
rect 8852 23060 8904 23112
rect 9588 23103 9640 23112
rect 9588 23069 9597 23103
rect 9597 23069 9631 23103
rect 9631 23069 9640 23103
rect 9588 23060 9640 23069
rect 8392 22992 8444 23044
rect 10232 22992 10284 23044
rect 15384 23137 15393 23171
rect 15393 23137 15427 23171
rect 15427 23137 15436 23171
rect 15384 23128 15436 23137
rect 15936 23128 15988 23180
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 17408 23128 17460 23180
rect 19340 23128 19392 23180
rect 20444 23128 20496 23180
rect 20904 23128 20956 23180
rect 21732 23128 21784 23180
rect 22192 23128 22244 23180
rect 15108 23060 15160 23112
rect 16396 23060 16448 23112
rect 16580 22992 16632 23044
rect 16764 23103 16816 23112
rect 16764 23069 16773 23103
rect 16773 23069 16807 23103
rect 16807 23069 16816 23103
rect 17500 23103 17552 23112
rect 16764 23060 16816 23069
rect 17500 23069 17509 23103
rect 17509 23069 17543 23103
rect 17543 23069 17552 23103
rect 17500 23060 17552 23069
rect 3424 22924 3476 22976
rect 4896 22924 4948 22976
rect 7840 22924 7892 22976
rect 9404 22924 9456 22976
rect 14464 22924 14516 22976
rect 15108 22924 15160 22976
rect 15844 22924 15896 22976
rect 16120 22924 16172 22976
rect 17132 22992 17184 23044
rect 19432 22992 19484 23044
rect 20260 22992 20312 23044
rect 21272 23103 21324 23112
rect 21272 23069 21281 23103
rect 21281 23069 21315 23103
rect 21315 23069 21324 23103
rect 21272 23060 21324 23069
rect 17960 22924 18012 22976
rect 20076 22924 20128 22976
rect 22376 23060 22428 23112
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 3700 22720 3752 22772
rect 5908 22720 5960 22772
rect 10232 22763 10284 22772
rect 10232 22729 10241 22763
rect 10241 22729 10275 22763
rect 10275 22729 10284 22763
rect 10232 22720 10284 22729
rect 15568 22763 15620 22772
rect 15568 22729 15577 22763
rect 15577 22729 15611 22763
rect 15611 22729 15620 22763
rect 15568 22720 15620 22729
rect 16580 22720 16632 22772
rect 16764 22720 16816 22772
rect 17132 22763 17184 22772
rect 17132 22729 17141 22763
rect 17141 22729 17175 22763
rect 17175 22729 17184 22763
rect 17132 22720 17184 22729
rect 17408 22720 17460 22772
rect 18972 22720 19024 22772
rect 20720 22720 20772 22772
rect 23480 22720 23532 22772
rect 3424 22695 3476 22704
rect 3424 22661 3433 22695
rect 3433 22661 3467 22695
rect 3467 22661 3476 22695
rect 3424 22652 3476 22661
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2964 22627 3016 22636
rect 2780 22584 2832 22593
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 3516 22584 3568 22636
rect 4344 22627 4396 22636
rect 4344 22593 4353 22627
rect 4353 22593 4387 22627
rect 4387 22593 4396 22627
rect 4344 22584 4396 22593
rect 4620 22584 4672 22636
rect 4804 22584 4856 22636
rect 5816 22652 5868 22704
rect 6552 22652 6604 22704
rect 6460 22584 6512 22636
rect 9496 22584 9548 22636
rect 11152 22652 11204 22704
rect 12256 22652 12308 22704
rect 4988 22516 5040 22568
rect 5448 22516 5500 22568
rect 2688 22448 2740 22500
rect 4160 22491 4212 22500
rect 2872 22423 2924 22432
rect 2872 22389 2881 22423
rect 2881 22389 2915 22423
rect 2915 22389 2924 22423
rect 2872 22380 2924 22389
rect 3332 22380 3384 22432
rect 4160 22457 4169 22491
rect 4169 22457 4203 22491
rect 4203 22457 4212 22491
rect 4160 22448 4212 22457
rect 4344 22380 4396 22432
rect 7840 22380 7892 22432
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 15660 22652 15712 22704
rect 17408 22627 17460 22636
rect 17408 22593 17417 22627
rect 17417 22593 17451 22627
rect 17451 22593 17460 22627
rect 17408 22584 17460 22593
rect 19248 22652 19300 22704
rect 20352 22652 20404 22704
rect 21272 22652 21324 22704
rect 21824 22652 21876 22704
rect 17592 22627 17644 22636
rect 17592 22593 17601 22627
rect 17601 22593 17635 22627
rect 17635 22593 17644 22627
rect 17592 22584 17644 22593
rect 12256 22559 12308 22568
rect 12256 22525 12265 22559
rect 12265 22525 12299 22559
rect 12299 22525 12308 22559
rect 12256 22516 12308 22525
rect 12716 22516 12768 22568
rect 15292 22516 15344 22568
rect 15844 22516 15896 22568
rect 18236 22584 18288 22636
rect 18604 22584 18656 22636
rect 19432 22627 19484 22636
rect 19432 22593 19441 22627
rect 19441 22593 19475 22627
rect 19475 22593 19484 22627
rect 19432 22584 19484 22593
rect 20260 22627 20312 22636
rect 20260 22593 20269 22627
rect 20269 22593 20303 22627
rect 20303 22593 20312 22627
rect 20260 22584 20312 22593
rect 19984 22516 20036 22568
rect 20444 22516 20496 22568
rect 20996 22559 21048 22568
rect 20996 22525 21005 22559
rect 21005 22525 21039 22559
rect 21039 22525 21048 22559
rect 20996 22516 21048 22525
rect 21640 22584 21692 22636
rect 21732 22516 21784 22568
rect 22192 22559 22244 22568
rect 22192 22525 22201 22559
rect 22201 22525 22235 22559
rect 22235 22525 22244 22559
rect 22192 22516 22244 22525
rect 10600 22491 10652 22500
rect 10600 22457 10609 22491
rect 10609 22457 10643 22491
rect 10643 22457 10652 22491
rect 10600 22448 10652 22457
rect 11152 22448 11204 22500
rect 11796 22491 11848 22500
rect 11796 22457 11805 22491
rect 11805 22457 11839 22491
rect 11839 22457 11848 22491
rect 11796 22448 11848 22457
rect 12808 22448 12860 22500
rect 14280 22448 14332 22500
rect 18696 22448 18748 22500
rect 11060 22380 11112 22432
rect 15752 22380 15804 22432
rect 21548 22380 21600 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2320 22176 2372 22228
rect 9588 22219 9640 22228
rect 2136 22015 2188 22024
rect 2136 21981 2145 22015
rect 2145 21981 2179 22015
rect 2179 21981 2188 22015
rect 2136 21972 2188 21981
rect 2688 21972 2740 22024
rect 2964 22015 3016 22024
rect 2964 21981 2973 22015
rect 2973 21981 3007 22015
rect 3007 21981 3016 22015
rect 2964 21972 3016 21981
rect 3516 22108 3568 22160
rect 9588 22185 9597 22219
rect 9597 22185 9631 22219
rect 9631 22185 9640 22219
rect 9588 22176 9640 22185
rect 12256 22176 12308 22228
rect 12716 22219 12768 22228
rect 12716 22185 12725 22219
rect 12725 22185 12759 22219
rect 12759 22185 12768 22219
rect 12716 22176 12768 22185
rect 21640 22176 21692 22228
rect 4068 22040 4120 22092
rect 3424 22015 3476 22024
rect 3424 21981 3433 22015
rect 3433 21981 3467 22015
rect 3467 21981 3476 22015
rect 4252 22015 4304 22024
rect 3424 21972 3476 21981
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 4896 22108 4948 22160
rect 6092 22108 6144 22160
rect 7840 22108 7892 22160
rect 8300 22151 8352 22160
rect 8300 22117 8309 22151
rect 8309 22117 8343 22151
rect 8343 22117 8352 22151
rect 8300 22108 8352 22117
rect 4896 22015 4948 22024
rect 4896 21981 4905 22015
rect 4905 21981 4939 22015
rect 4939 21981 4948 22015
rect 4896 21972 4948 21981
rect 5448 21972 5500 22024
rect 8944 22040 8996 22092
rect 11060 22040 11112 22092
rect 12348 22083 12400 22092
rect 12348 22049 12357 22083
rect 12357 22049 12391 22083
rect 12391 22049 12400 22083
rect 12348 22040 12400 22049
rect 17500 22108 17552 22160
rect 9588 21972 9640 22024
rect 10692 21972 10744 22024
rect 11244 21972 11296 22024
rect 12440 22015 12492 22024
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12440 21972 12492 21981
rect 12624 21972 12676 22024
rect 13636 22015 13688 22024
rect 13636 21981 13645 22015
rect 13645 21981 13679 22015
rect 13679 21981 13688 22015
rect 13636 21972 13688 21981
rect 14280 22015 14332 22024
rect 3608 21904 3660 21956
rect 5632 21904 5684 21956
rect 3240 21836 3292 21888
rect 6644 21836 6696 21888
rect 9404 21904 9456 21956
rect 11060 21904 11112 21956
rect 11888 21904 11940 21956
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 17224 22040 17276 22092
rect 17868 22040 17920 22092
rect 15384 21972 15436 22024
rect 16488 21972 16540 22024
rect 17040 21972 17092 22024
rect 17592 21972 17644 22024
rect 18512 21972 18564 22024
rect 18696 22015 18748 22024
rect 18696 21981 18705 22015
rect 18705 21981 18739 22015
rect 18739 21981 18748 22015
rect 18696 21972 18748 21981
rect 19984 21972 20036 22024
rect 21548 22015 21600 22024
rect 21548 21981 21557 22015
rect 21557 21981 21591 22015
rect 21591 21981 21600 22015
rect 21548 21972 21600 21981
rect 21732 22015 21784 22024
rect 21732 21981 21741 22015
rect 21741 21981 21775 22015
rect 21775 21981 21784 22015
rect 21732 21972 21784 21981
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 23204 21972 23256 22024
rect 13912 21904 13964 21956
rect 15752 21904 15804 21956
rect 15936 21904 15988 21956
rect 9864 21836 9916 21888
rect 11336 21879 11388 21888
rect 11336 21845 11345 21879
rect 11345 21845 11379 21879
rect 11379 21845 11388 21879
rect 11336 21836 11388 21845
rect 15200 21836 15252 21888
rect 17040 21836 17092 21888
rect 17408 21836 17460 21888
rect 20168 21836 20220 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2780 21675 2832 21684
rect 2780 21641 2789 21675
rect 2789 21641 2823 21675
rect 2823 21641 2832 21675
rect 2780 21632 2832 21641
rect 4252 21632 4304 21684
rect 7380 21675 7432 21684
rect 7380 21641 7389 21675
rect 7389 21641 7423 21675
rect 7423 21641 7432 21675
rect 7380 21632 7432 21641
rect 2136 21564 2188 21616
rect 2872 21496 2924 21548
rect 3056 21428 3108 21480
rect 3332 21471 3384 21480
rect 3332 21437 3341 21471
rect 3341 21437 3375 21471
rect 3375 21437 3384 21471
rect 3332 21428 3384 21437
rect 4712 21496 4764 21548
rect 4988 21564 5040 21616
rect 9588 21632 9640 21684
rect 9864 21632 9916 21684
rect 12532 21632 12584 21684
rect 13636 21632 13688 21684
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 11980 21564 12032 21616
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 8392 21539 8444 21548
rect 8392 21505 8401 21539
rect 8401 21505 8435 21539
rect 8435 21505 8444 21539
rect 8392 21496 8444 21505
rect 8576 21539 8628 21548
rect 8576 21505 8585 21539
rect 8585 21505 8619 21539
rect 8619 21505 8628 21539
rect 8576 21496 8628 21505
rect 8668 21539 8720 21548
rect 8668 21505 8677 21539
rect 8677 21505 8711 21539
rect 8711 21505 8720 21539
rect 8852 21539 8904 21548
rect 8668 21496 8720 21505
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 8944 21539 8996 21548
rect 8944 21505 8953 21539
rect 8953 21505 8987 21539
rect 8987 21505 8996 21539
rect 8944 21496 8996 21505
rect 9864 21496 9916 21548
rect 10876 21496 10928 21548
rect 11796 21496 11848 21548
rect 15476 21564 15528 21616
rect 15660 21632 15712 21684
rect 17408 21632 17460 21684
rect 17868 21632 17920 21684
rect 22008 21632 22060 21684
rect 23204 21632 23256 21684
rect 19432 21564 19484 21616
rect 15200 21539 15252 21548
rect 15200 21505 15209 21539
rect 15209 21505 15243 21539
rect 15243 21505 15252 21539
rect 15200 21496 15252 21505
rect 16948 21496 17000 21548
rect 17684 21496 17736 21548
rect 20168 21564 20220 21616
rect 20904 21564 20956 21616
rect 21732 21564 21784 21616
rect 19616 21539 19668 21548
rect 19616 21505 19625 21539
rect 19625 21505 19659 21539
rect 19659 21505 19668 21539
rect 19616 21496 19668 21505
rect 20536 21496 20588 21548
rect 21824 21496 21876 21548
rect 23020 21496 23072 21548
rect 4804 21471 4856 21480
rect 4804 21437 4813 21471
rect 4813 21437 4847 21471
rect 4847 21437 4856 21471
rect 4804 21428 4856 21437
rect 6092 21428 6144 21480
rect 6000 21403 6052 21412
rect 6000 21369 6009 21403
rect 6009 21369 6043 21403
rect 6043 21369 6052 21403
rect 6000 21360 6052 21369
rect 7380 21428 7432 21480
rect 9312 21428 9364 21480
rect 10784 21471 10836 21480
rect 10784 21437 10793 21471
rect 10793 21437 10827 21471
rect 10827 21437 10836 21471
rect 10784 21428 10836 21437
rect 7932 21360 7984 21412
rect 8852 21360 8904 21412
rect 8484 21292 8536 21344
rect 12532 21428 12584 21480
rect 17040 21428 17092 21480
rect 19984 21428 20036 21480
rect 22192 21428 22244 21480
rect 11336 21360 11388 21412
rect 11152 21335 11204 21344
rect 11152 21301 11161 21335
rect 11161 21301 11195 21335
rect 11195 21301 11204 21335
rect 11152 21292 11204 21301
rect 15292 21335 15344 21344
rect 15292 21301 15301 21335
rect 15301 21301 15335 21335
rect 15335 21301 15344 21335
rect 15292 21292 15344 21301
rect 15384 21335 15436 21344
rect 15384 21301 15393 21335
rect 15393 21301 15427 21335
rect 15427 21301 15436 21335
rect 15384 21292 15436 21301
rect 16764 21292 16816 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6736 21088 6788 21140
rect 7104 21131 7156 21140
rect 6276 21020 6328 21072
rect 7104 21097 7113 21131
rect 7113 21097 7147 21131
rect 7147 21097 7156 21131
rect 7104 21088 7156 21097
rect 7932 21131 7984 21140
rect 7932 21097 7941 21131
rect 7941 21097 7975 21131
rect 7975 21097 7984 21131
rect 7932 21088 7984 21097
rect 7012 21020 7064 21072
rect 8576 21088 8628 21140
rect 9404 21088 9456 21140
rect 10600 21088 10652 21140
rect 11152 21088 11204 21140
rect 4252 20952 4304 21004
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 3976 20884 4028 20936
rect 5632 20884 5684 20936
rect 5908 20927 5960 20936
rect 5908 20893 5917 20927
rect 5917 20893 5951 20927
rect 5951 20893 5960 20927
rect 5908 20884 5960 20893
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6000 20884 6052 20893
rect 6368 20884 6420 20936
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 6552 20884 6604 20893
rect 6920 20884 6972 20936
rect 8300 21020 8352 21072
rect 12256 21088 12308 21140
rect 12440 21088 12492 21140
rect 7840 20952 7892 21004
rect 9680 20952 9732 21004
rect 11520 20952 11572 21004
rect 15292 21088 15344 21140
rect 15844 21088 15896 21140
rect 17684 21131 17736 21140
rect 17684 21097 17693 21131
rect 17693 21097 17727 21131
rect 17727 21097 17736 21131
rect 17684 21088 17736 21097
rect 18696 21088 18748 21140
rect 20996 21088 21048 21140
rect 21272 21088 21324 21140
rect 23020 21131 23072 21140
rect 23020 21097 23029 21131
rect 23029 21097 23063 21131
rect 23063 21097 23072 21131
rect 23020 21088 23072 21097
rect 17500 21020 17552 21072
rect 11888 20995 11940 21004
rect 11888 20961 11897 20995
rect 11897 20961 11931 20995
rect 11931 20961 11940 20995
rect 11888 20952 11940 20961
rect 2964 20816 3016 20868
rect 6092 20816 6144 20868
rect 8484 20884 8536 20936
rect 10600 20884 10652 20936
rect 10968 20927 11020 20936
rect 10968 20893 10977 20927
rect 10977 20893 11011 20927
rect 11011 20893 11020 20927
rect 10968 20884 11020 20893
rect 11244 20884 11296 20936
rect 8668 20816 8720 20868
rect 9680 20816 9732 20868
rect 11060 20816 11112 20868
rect 11704 20927 11756 20936
rect 11704 20893 11713 20927
rect 11713 20893 11747 20927
rect 11747 20893 11756 20927
rect 12348 20927 12400 20936
rect 11704 20884 11756 20893
rect 12348 20893 12357 20927
rect 12357 20893 12391 20927
rect 12391 20893 12400 20927
rect 12348 20884 12400 20893
rect 12532 20927 12584 20936
rect 12532 20893 12541 20927
rect 12541 20893 12575 20927
rect 12575 20893 12584 20927
rect 12532 20884 12584 20893
rect 14648 20952 14700 21004
rect 16764 20952 16816 21004
rect 15660 20884 15712 20936
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 18512 21020 18564 21072
rect 19616 21063 19668 21072
rect 19616 21029 19625 21063
rect 19625 21029 19659 21063
rect 19659 21029 19668 21063
rect 19616 21020 19668 21029
rect 15936 20816 15988 20868
rect 17868 20884 17920 20936
rect 18972 20952 19024 21004
rect 20260 21020 20312 21072
rect 22192 21020 22244 21072
rect 20444 20952 20496 21004
rect 21732 20952 21784 21004
rect 18328 20884 18380 20936
rect 19248 20884 19300 20936
rect 20168 20884 20220 20936
rect 20352 20884 20404 20936
rect 20904 20884 20956 20936
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 21088 20884 21140 20893
rect 1768 20791 1820 20800
rect 1768 20757 1777 20791
rect 1777 20757 1811 20791
rect 1811 20757 1820 20791
rect 1768 20748 1820 20757
rect 3424 20791 3476 20800
rect 3424 20757 3433 20791
rect 3433 20757 3467 20791
rect 3467 20757 3476 20791
rect 3424 20748 3476 20757
rect 7012 20748 7064 20800
rect 9772 20748 9824 20800
rect 12164 20748 12216 20800
rect 15108 20748 15160 20800
rect 17592 20816 17644 20868
rect 17500 20748 17552 20800
rect 18328 20748 18380 20800
rect 21456 20791 21508 20800
rect 21456 20757 21465 20791
rect 21465 20757 21499 20791
rect 21499 20757 21508 20791
rect 21456 20748 21508 20757
rect 22928 20748 22980 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5908 20544 5960 20596
rect 6460 20544 6512 20596
rect 8576 20544 8628 20596
rect 9588 20544 9640 20596
rect 10784 20544 10836 20596
rect 11520 20544 11572 20596
rect 13176 20544 13228 20596
rect 14740 20544 14792 20596
rect 15936 20544 15988 20596
rect 18696 20544 18748 20596
rect 3056 20476 3108 20528
rect 2228 20408 2280 20460
rect 2320 20451 2372 20460
rect 2320 20417 2329 20451
rect 2329 20417 2363 20451
rect 2363 20417 2372 20451
rect 5448 20476 5500 20528
rect 2320 20408 2372 20417
rect 3884 20408 3936 20460
rect 4252 20451 4304 20460
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 4252 20408 4304 20417
rect 4620 20408 4672 20460
rect 5264 20408 5316 20460
rect 3424 20383 3476 20392
rect 3424 20349 3433 20383
rect 3433 20349 3467 20383
rect 3467 20349 3476 20383
rect 3424 20340 3476 20349
rect 3976 20340 4028 20392
rect 6092 20408 6144 20460
rect 8484 20476 8536 20528
rect 11796 20476 11848 20528
rect 7380 20451 7432 20460
rect 7380 20417 7389 20451
rect 7389 20417 7423 20451
rect 7423 20417 7432 20451
rect 7380 20408 7432 20417
rect 8300 20408 8352 20460
rect 9312 20408 9364 20460
rect 11060 20408 11112 20460
rect 11704 20408 11756 20460
rect 11980 20408 12032 20460
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 14280 20408 14332 20460
rect 15844 20476 15896 20528
rect 14832 20408 14884 20460
rect 15660 20408 15712 20460
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 16304 20451 16356 20460
rect 16304 20417 16313 20451
rect 16313 20417 16347 20451
rect 16347 20417 16356 20451
rect 17776 20451 17828 20460
rect 16304 20408 16356 20417
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 21456 20544 21508 20596
rect 6828 20340 6880 20392
rect 7472 20340 7524 20392
rect 10692 20340 10744 20392
rect 13176 20340 13228 20392
rect 14464 20383 14516 20392
rect 14464 20349 14473 20383
rect 14473 20349 14507 20383
rect 14507 20349 14516 20383
rect 14464 20340 14516 20349
rect 14648 20383 14700 20392
rect 14648 20349 14657 20383
rect 14657 20349 14691 20383
rect 14691 20349 14700 20383
rect 14648 20340 14700 20349
rect 3056 20272 3108 20324
rect 6092 20272 6144 20324
rect 9864 20315 9916 20324
rect 9864 20281 9873 20315
rect 9873 20281 9907 20315
rect 9907 20281 9916 20315
rect 9864 20272 9916 20281
rect 10968 20272 11020 20324
rect 11888 20272 11940 20324
rect 11980 20315 12032 20324
rect 11980 20281 11989 20315
rect 11989 20281 12023 20315
rect 12023 20281 12032 20315
rect 11980 20272 12032 20281
rect 14924 20272 14976 20324
rect 16304 20272 16356 20324
rect 18052 20272 18104 20324
rect 18144 20272 18196 20324
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 2136 20247 2188 20256
rect 2136 20213 2145 20247
rect 2145 20213 2179 20247
rect 2179 20213 2188 20247
rect 2136 20204 2188 20213
rect 3240 20247 3292 20256
rect 3240 20213 3249 20247
rect 3249 20213 3283 20247
rect 3283 20213 3292 20247
rect 3240 20204 3292 20213
rect 4068 20204 4120 20256
rect 5632 20204 5684 20256
rect 9680 20247 9732 20256
rect 9680 20213 9689 20247
rect 9689 20213 9723 20247
rect 9723 20213 9732 20247
rect 9680 20204 9732 20213
rect 11060 20247 11112 20256
rect 11060 20213 11069 20247
rect 11069 20213 11103 20247
rect 11103 20213 11112 20247
rect 11060 20204 11112 20213
rect 13084 20204 13136 20256
rect 14556 20204 14608 20256
rect 15660 20204 15712 20256
rect 15844 20204 15896 20256
rect 17868 20204 17920 20256
rect 18604 20247 18656 20256
rect 18604 20213 18613 20247
rect 18613 20213 18647 20247
rect 18647 20213 18656 20247
rect 18604 20204 18656 20213
rect 19432 20204 19484 20256
rect 20168 20247 20220 20256
rect 20168 20213 20177 20247
rect 20177 20213 20211 20247
rect 20211 20213 20220 20247
rect 20168 20204 20220 20213
rect 20352 20247 20404 20256
rect 20352 20213 20361 20247
rect 20361 20213 20395 20247
rect 20395 20213 20404 20247
rect 20352 20204 20404 20213
rect 20536 20408 20588 20460
rect 20996 20451 21048 20460
rect 20996 20417 21005 20451
rect 21005 20417 21039 20451
rect 21039 20417 21048 20451
rect 20996 20408 21048 20417
rect 21364 20408 21416 20460
rect 22928 20451 22980 20460
rect 20904 20340 20956 20392
rect 21272 20272 21324 20324
rect 22928 20417 22937 20451
rect 22937 20417 22971 20451
rect 22971 20417 22980 20451
rect 22928 20408 22980 20417
rect 22100 20204 22152 20256
rect 22744 20247 22796 20256
rect 22744 20213 22753 20247
rect 22753 20213 22787 20247
rect 22787 20213 22796 20247
rect 22744 20204 22796 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2228 20000 2280 20052
rect 4804 20000 4856 20052
rect 6276 20000 6328 20052
rect 6552 20000 6604 20052
rect 7380 20000 7432 20052
rect 2964 19975 3016 19984
rect 2964 19941 2973 19975
rect 2973 19941 3007 19975
rect 3007 19941 3016 19975
rect 2964 19932 3016 19941
rect 3240 19864 3292 19916
rect 6460 19907 6512 19916
rect 2136 19796 2188 19848
rect 3424 19796 3476 19848
rect 6460 19873 6469 19907
rect 6469 19873 6503 19907
rect 6503 19873 6512 19907
rect 6460 19864 6512 19873
rect 6368 19839 6420 19848
rect 4896 19728 4948 19780
rect 1860 19660 1912 19712
rect 4068 19660 4120 19712
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 6552 19796 6604 19848
rect 7656 19864 7708 19916
rect 11060 20000 11112 20052
rect 15752 20000 15804 20052
rect 8484 19975 8536 19984
rect 8484 19941 8493 19975
rect 8493 19941 8527 19975
rect 8527 19941 8536 19975
rect 8484 19932 8536 19941
rect 10600 19932 10652 19984
rect 9588 19864 9640 19916
rect 11888 19932 11940 19984
rect 14924 19975 14976 19984
rect 14924 19941 14933 19975
rect 14933 19941 14967 19975
rect 14967 19941 14976 19975
rect 14924 19932 14976 19941
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 5724 19728 5776 19780
rect 7748 19728 7800 19780
rect 11796 19796 11848 19848
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 12072 19796 12124 19848
rect 12716 19796 12768 19848
rect 14740 19864 14792 19916
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 13268 19839 13320 19848
rect 13268 19805 13275 19839
rect 13275 19805 13320 19839
rect 13268 19796 13320 19805
rect 13728 19796 13780 19848
rect 9404 19728 9456 19780
rect 13360 19771 13412 19780
rect 13360 19737 13369 19771
rect 13369 19737 13403 19771
rect 13403 19737 13412 19771
rect 13360 19728 13412 19737
rect 13820 19728 13872 19780
rect 18144 20000 18196 20052
rect 18328 20043 18380 20052
rect 18328 20009 18337 20043
rect 18337 20009 18371 20043
rect 18371 20009 18380 20043
rect 18328 20000 18380 20009
rect 20352 20000 20404 20052
rect 21088 20000 21140 20052
rect 21364 20000 21416 20052
rect 16304 19932 16356 19984
rect 20076 19975 20128 19984
rect 20076 19941 20085 19975
rect 20085 19941 20119 19975
rect 20119 19941 20128 19975
rect 20076 19932 20128 19941
rect 15936 19864 15988 19916
rect 15200 19796 15252 19848
rect 16028 19796 16080 19848
rect 16764 19864 16816 19916
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 18604 19864 18656 19916
rect 20536 19864 20588 19916
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 14280 19660 14332 19712
rect 17684 19728 17736 19780
rect 17868 19728 17920 19780
rect 16212 19660 16264 19712
rect 16304 19660 16356 19712
rect 18420 19660 18472 19712
rect 19340 19728 19392 19780
rect 20628 19796 20680 19848
rect 20996 19796 21048 19848
rect 21180 19796 21232 19848
rect 22744 19796 22796 19848
rect 21272 19660 21324 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3976 19456 4028 19508
rect 1952 19388 2004 19440
rect 5448 19456 5500 19508
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 4712 19388 4764 19440
rect 6000 19388 6052 19440
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 5632 19320 5684 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 6644 19320 6696 19372
rect 8300 19456 8352 19508
rect 13268 19456 13320 19508
rect 14832 19499 14884 19508
rect 7564 19388 7616 19440
rect 12716 19388 12768 19440
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 15660 19456 15712 19508
rect 15752 19456 15804 19508
rect 16120 19456 16172 19508
rect 18052 19499 18104 19508
rect 2964 19252 3016 19304
rect 5448 19252 5500 19304
rect 1860 19227 1912 19236
rect 1860 19193 1869 19227
rect 1869 19193 1903 19227
rect 1903 19193 1912 19227
rect 1860 19184 1912 19193
rect 5540 19184 5592 19236
rect 4620 19116 4672 19168
rect 6736 19116 6788 19168
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 7288 19252 7340 19304
rect 8852 19295 8904 19304
rect 8852 19261 8861 19295
rect 8861 19261 8895 19295
rect 8895 19261 8904 19295
rect 8852 19252 8904 19261
rect 9404 19295 9456 19304
rect 9404 19261 9413 19295
rect 9413 19261 9447 19295
rect 9447 19261 9456 19295
rect 9404 19252 9456 19261
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 12808 19363 12860 19372
rect 11060 19320 11112 19329
rect 12808 19329 12817 19363
rect 12817 19329 12851 19363
rect 12851 19329 12860 19363
rect 12808 19320 12860 19329
rect 13268 19363 13320 19372
rect 13268 19329 13277 19363
rect 13277 19329 13311 19363
rect 13311 19329 13320 19363
rect 13268 19320 13320 19329
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 15844 19388 15896 19440
rect 13820 19363 13872 19372
rect 13820 19329 13829 19363
rect 13829 19329 13863 19363
rect 13863 19329 13872 19363
rect 13820 19320 13872 19329
rect 14464 19320 14516 19372
rect 11244 19252 11296 19304
rect 13728 19295 13780 19304
rect 13728 19261 13737 19295
rect 13737 19261 13771 19295
rect 13771 19261 13780 19295
rect 13728 19252 13780 19261
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 10876 19227 10928 19236
rect 10876 19193 10885 19227
rect 10885 19193 10919 19227
rect 10919 19193 10928 19227
rect 10876 19184 10928 19193
rect 18052 19465 18061 19499
rect 18061 19465 18095 19499
rect 18095 19465 18104 19499
rect 18052 19456 18104 19465
rect 18144 19456 18196 19508
rect 20260 19456 20312 19508
rect 20168 19388 20220 19440
rect 20628 19388 20680 19440
rect 17776 19320 17828 19372
rect 18144 19363 18196 19372
rect 18144 19329 18153 19363
rect 18153 19329 18187 19363
rect 18187 19329 18196 19363
rect 18696 19363 18748 19372
rect 18144 19320 18196 19329
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 19340 19320 19392 19372
rect 17592 19252 17644 19304
rect 17868 19252 17920 19304
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 20996 19320 21048 19372
rect 21364 19320 21416 19372
rect 22100 19320 22152 19372
rect 21088 19252 21140 19304
rect 7932 19159 7984 19168
rect 7932 19125 7941 19159
rect 7941 19125 7975 19159
rect 7975 19125 7984 19159
rect 7932 19116 7984 19125
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 11152 19116 11204 19168
rect 12624 19159 12676 19168
rect 12624 19125 12633 19159
rect 12633 19125 12667 19159
rect 12667 19125 12676 19159
rect 12624 19116 12676 19125
rect 13636 19159 13688 19168
rect 13636 19125 13645 19159
rect 13645 19125 13679 19159
rect 13679 19125 13688 19159
rect 13636 19116 13688 19125
rect 13912 19116 13964 19168
rect 17316 19116 17368 19168
rect 17960 19116 18012 19168
rect 18972 19116 19024 19168
rect 20352 19116 20404 19168
rect 20536 19159 20588 19168
rect 20536 19125 20545 19159
rect 20545 19125 20579 19159
rect 20579 19125 20588 19159
rect 20536 19116 20588 19125
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 38292 19159 38344 19168
rect 38292 19125 38301 19159
rect 38301 19125 38335 19159
rect 38335 19125 38344 19159
rect 38292 19116 38344 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3240 18912 3292 18964
rect 5632 18955 5684 18964
rect 5632 18921 5641 18955
rect 5641 18921 5675 18955
rect 5675 18921 5684 18955
rect 5632 18912 5684 18921
rect 6920 18912 6972 18964
rect 8300 18912 8352 18964
rect 8852 18912 8904 18964
rect 13636 18912 13688 18964
rect 15476 18912 15528 18964
rect 11244 18844 11296 18896
rect 12440 18844 12492 18896
rect 16948 18912 17000 18964
rect 17684 18955 17736 18964
rect 17684 18921 17693 18955
rect 17693 18921 17727 18955
rect 17727 18921 17736 18955
rect 17684 18912 17736 18921
rect 17776 18912 17828 18964
rect 19340 18912 19392 18964
rect 21364 18912 21416 18964
rect 16304 18844 16356 18896
rect 16580 18844 16632 18896
rect 18144 18844 18196 18896
rect 19248 18844 19300 18896
rect 3056 18776 3108 18828
rect 2964 18708 3016 18760
rect 4436 18751 4488 18760
rect 4436 18717 4445 18751
rect 4445 18717 4479 18751
rect 4479 18717 4488 18751
rect 4436 18708 4488 18717
rect 6644 18776 6696 18828
rect 7472 18819 7524 18828
rect 7472 18785 7481 18819
rect 7481 18785 7515 18819
rect 7515 18785 7524 18819
rect 7472 18776 7524 18785
rect 7932 18776 7984 18828
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 5908 18640 5960 18692
rect 4620 18572 4672 18624
rect 7656 18708 7708 18760
rect 7748 18708 7800 18760
rect 8116 18708 8168 18760
rect 15292 18776 15344 18828
rect 16396 18776 16448 18828
rect 12900 18708 12952 18760
rect 14096 18708 14148 18760
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 17776 18708 17828 18760
rect 17960 18708 18012 18760
rect 18144 18751 18196 18760
rect 18144 18717 18153 18751
rect 18153 18717 18187 18751
rect 18187 18717 18196 18751
rect 18144 18708 18196 18717
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 20168 18751 20220 18760
rect 20168 18717 20177 18751
rect 20177 18717 20211 18751
rect 20211 18717 20220 18751
rect 20168 18708 20220 18717
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 21180 18751 21232 18760
rect 21180 18717 21189 18751
rect 21189 18717 21223 18751
rect 21223 18717 21232 18751
rect 21180 18708 21232 18717
rect 22008 18708 22060 18760
rect 10784 18640 10836 18692
rect 13636 18640 13688 18692
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 7104 18572 7156 18581
rect 7564 18572 7616 18624
rect 7840 18572 7892 18624
rect 9956 18572 10008 18624
rect 12164 18572 12216 18624
rect 14004 18640 14056 18692
rect 14280 18683 14332 18692
rect 14280 18649 14289 18683
rect 14289 18649 14323 18683
rect 14323 18649 14332 18683
rect 14280 18640 14332 18649
rect 17500 18640 17552 18692
rect 17592 18640 17644 18692
rect 20720 18640 20772 18692
rect 13912 18572 13964 18624
rect 16488 18572 16540 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17132 18572 17184 18581
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4712 18368 4764 18420
rect 6276 18368 6328 18420
rect 8116 18368 8168 18420
rect 10784 18411 10836 18420
rect 10784 18377 10793 18411
rect 10793 18377 10827 18411
rect 10827 18377 10836 18411
rect 10784 18368 10836 18377
rect 4436 18232 4488 18284
rect 4620 18275 4672 18284
rect 4620 18241 4629 18275
rect 4629 18241 4663 18275
rect 4663 18241 4672 18275
rect 4620 18232 4672 18241
rect 6092 18300 6144 18352
rect 6644 18300 6696 18352
rect 7104 18300 7156 18352
rect 8392 18300 8444 18352
rect 10692 18343 10744 18352
rect 10692 18309 10701 18343
rect 10701 18309 10735 18343
rect 10735 18309 10744 18343
rect 10692 18300 10744 18309
rect 12992 18300 13044 18352
rect 5540 18275 5592 18284
rect 5540 18241 5549 18275
rect 5549 18241 5583 18275
rect 5583 18241 5592 18275
rect 5540 18232 5592 18241
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8024 18275 8076 18284
rect 8024 18241 8033 18275
rect 8033 18241 8067 18275
rect 8067 18241 8076 18275
rect 8024 18232 8076 18241
rect 8484 18232 8536 18284
rect 11888 18275 11940 18284
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 12716 18232 12768 18284
rect 3056 18207 3108 18216
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 3056 18164 3108 18173
rect 5724 18164 5776 18216
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 8208 18164 8260 18216
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 3884 18096 3936 18148
rect 13912 18368 13964 18420
rect 14096 18411 14148 18420
rect 14096 18377 14105 18411
rect 14105 18377 14139 18411
rect 14139 18377 14148 18411
rect 14096 18368 14148 18377
rect 18328 18368 18380 18420
rect 20444 18368 20496 18420
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 15568 18300 15620 18352
rect 17776 18343 17828 18352
rect 17776 18309 17785 18343
rect 17785 18309 17819 18343
rect 17819 18309 17828 18343
rect 17776 18300 17828 18309
rect 19064 18300 19116 18352
rect 20260 18300 20312 18352
rect 13544 18275 13596 18284
rect 13544 18241 13554 18275
rect 13554 18241 13588 18275
rect 13588 18241 13596 18275
rect 13544 18232 13596 18241
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 14004 18232 14056 18284
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 17500 18232 17552 18284
rect 18604 18232 18656 18284
rect 19984 18232 20036 18284
rect 4804 18028 4856 18080
rect 6736 18071 6788 18080
rect 6736 18037 6745 18071
rect 6745 18037 6779 18071
rect 6779 18037 6788 18071
rect 6736 18028 6788 18037
rect 7840 18028 7892 18080
rect 14096 18164 14148 18216
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 15384 18164 15436 18216
rect 17960 18096 18012 18148
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 12532 18028 12584 18080
rect 12992 18071 13044 18080
rect 12992 18037 13001 18071
rect 13001 18037 13035 18071
rect 13035 18037 13044 18071
rect 12992 18028 13044 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4620 17824 4672 17876
rect 7932 17824 7984 17876
rect 12532 17824 12584 17876
rect 12808 17824 12860 17876
rect 13268 17824 13320 17876
rect 6644 17756 6696 17808
rect 10692 17756 10744 17808
rect 13728 17824 13780 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15476 17824 15528 17876
rect 17776 17824 17828 17876
rect 17960 17867 18012 17876
rect 17960 17833 17969 17867
rect 17969 17833 18003 17867
rect 18003 17833 18012 17867
rect 17960 17824 18012 17833
rect 18144 17824 18196 17876
rect 5540 17688 5592 17740
rect 8116 17688 8168 17740
rect 13636 17756 13688 17808
rect 14464 17756 14516 17808
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 4712 17620 4764 17672
rect 4804 17620 4856 17672
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 5264 17620 5316 17672
rect 6736 17620 6788 17672
rect 7104 17620 7156 17672
rect 3148 17552 3200 17604
rect 7656 17620 7708 17672
rect 10600 17620 10652 17672
rect 12072 17620 12124 17672
rect 13176 17620 13228 17672
rect 14096 17688 14148 17740
rect 16856 17688 16908 17740
rect 13544 17620 13596 17672
rect 13820 17620 13872 17672
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 15292 17620 15344 17672
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 18236 17756 18288 17808
rect 16304 17620 16356 17629
rect 15476 17552 15528 17604
rect 18420 17595 18472 17604
rect 5356 17527 5408 17536
rect 5356 17493 5365 17527
rect 5365 17493 5399 17527
rect 5399 17493 5408 17527
rect 5356 17484 5408 17493
rect 7472 17484 7524 17536
rect 10416 17527 10468 17536
rect 10416 17493 10425 17527
rect 10425 17493 10459 17527
rect 10459 17493 10468 17527
rect 10416 17484 10468 17493
rect 10508 17484 10560 17536
rect 11704 17484 11756 17536
rect 12992 17484 13044 17536
rect 15660 17484 15712 17536
rect 18420 17561 18429 17595
rect 18429 17561 18463 17595
rect 18463 17561 18472 17595
rect 18420 17552 18472 17561
rect 18788 17527 18840 17536
rect 18788 17493 18797 17527
rect 18797 17493 18831 17527
rect 18831 17493 18840 17527
rect 18788 17484 18840 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 5540 17280 5592 17332
rect 7104 17323 7156 17332
rect 7104 17289 7113 17323
rect 7113 17289 7147 17323
rect 7147 17289 7156 17323
rect 7104 17280 7156 17289
rect 9772 17280 9824 17332
rect 1860 17076 1912 17128
rect 4068 17144 4120 17196
rect 5172 17212 5224 17264
rect 8392 17212 8444 17264
rect 9128 17212 9180 17264
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 7840 17187 7892 17196
rect 6736 17144 6788 17153
rect 7840 17153 7849 17187
rect 7849 17153 7883 17187
rect 7883 17153 7892 17187
rect 7840 17144 7892 17153
rect 10508 17212 10560 17264
rect 12624 17280 12676 17332
rect 12716 17280 12768 17332
rect 15016 17280 15068 17332
rect 16120 17280 16172 17332
rect 18420 17280 18472 17332
rect 11152 17212 11204 17264
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 14464 17187 14516 17196
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 11060 17076 11112 17128
rect 11888 17076 11940 17128
rect 15016 17144 15068 17196
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 15660 17144 15712 17196
rect 15752 17144 15804 17196
rect 16672 17144 16724 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 18328 17144 18380 17196
rect 16856 17076 16908 17128
rect 18420 17076 18472 17128
rect 9036 17008 9088 17060
rect 15108 17008 15160 17060
rect 18144 17008 18196 17060
rect 7380 16940 7432 16992
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 12808 16940 12860 16992
rect 13636 16940 13688 16992
rect 15936 16940 15988 16992
rect 16028 16940 16080 16992
rect 19248 16940 19300 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4068 16779 4120 16788
rect 4068 16745 4077 16779
rect 4077 16745 4111 16779
rect 4111 16745 4120 16779
rect 4068 16736 4120 16745
rect 6828 16736 6880 16788
rect 9404 16736 9456 16788
rect 11152 16779 11204 16788
rect 11152 16745 11161 16779
rect 11161 16745 11195 16779
rect 11195 16745 11204 16779
rect 11152 16736 11204 16745
rect 15292 16736 15344 16788
rect 16120 16736 16172 16788
rect 18328 16779 18380 16788
rect 18328 16745 18337 16779
rect 18337 16745 18371 16779
rect 18371 16745 18380 16779
rect 18328 16736 18380 16745
rect 9128 16643 9180 16652
rect 5356 16532 5408 16584
rect 6000 16532 6052 16584
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 15200 16668 15252 16720
rect 11888 16600 11940 16652
rect 12164 16600 12216 16652
rect 15568 16643 15620 16652
rect 8208 16532 8260 16584
rect 9956 16532 10008 16584
rect 7288 16507 7340 16516
rect 7288 16473 7322 16507
rect 7322 16473 7340 16507
rect 7288 16464 7340 16473
rect 12716 16532 12768 16584
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 18512 16668 18564 16720
rect 19064 16668 19116 16720
rect 11796 16464 11848 16516
rect 13544 16464 13596 16516
rect 15476 16464 15528 16516
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 16396 16575 16448 16584
rect 15752 16532 15804 16541
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 16488 16532 16540 16584
rect 17224 16532 17276 16584
rect 18052 16600 18104 16652
rect 18788 16532 18840 16584
rect 10968 16396 11020 16448
rect 12256 16396 12308 16448
rect 15660 16396 15712 16448
rect 17592 16464 17644 16516
rect 17316 16396 17368 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 7288 16192 7340 16244
rect 10784 16192 10836 16244
rect 11520 16192 11572 16244
rect 15384 16192 15436 16244
rect 15568 16192 15620 16244
rect 16304 16192 16356 16244
rect 10968 16167 11020 16176
rect 10968 16133 10977 16167
rect 10977 16133 11011 16167
rect 11011 16133 11020 16167
rect 10968 16124 11020 16133
rect 12624 16124 12676 16176
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 8760 16056 8812 16108
rect 10324 16056 10376 16108
rect 10876 16056 10928 16108
rect 11704 16056 11756 16108
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 15476 16124 15528 16176
rect 16488 16124 16540 16176
rect 12900 16056 12952 16108
rect 15108 16099 15160 16108
rect 15108 16065 15117 16099
rect 15117 16065 15151 16099
rect 15151 16065 15160 16099
rect 15108 16056 15160 16065
rect 15292 16099 15344 16108
rect 15292 16065 15301 16099
rect 15301 16065 15335 16099
rect 15335 16065 15344 16099
rect 15292 16056 15344 16065
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 17040 16167 17092 16176
rect 17040 16133 17065 16167
rect 17065 16133 17092 16167
rect 17592 16192 17644 16244
rect 19064 16235 19116 16244
rect 19064 16201 19073 16235
rect 19073 16201 19107 16235
rect 19107 16201 19116 16235
rect 19064 16192 19116 16201
rect 17040 16124 17092 16133
rect 17224 16056 17276 16108
rect 17408 16124 17460 16176
rect 18420 16124 18472 16176
rect 18512 16124 18564 16176
rect 22284 16124 22336 16176
rect 13544 16031 13596 16040
rect 10324 15920 10376 15972
rect 11336 15920 11388 15972
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 15384 16031 15436 16040
rect 15384 15997 15393 16031
rect 15393 15997 15427 16031
rect 15427 15997 15436 16031
rect 15384 15988 15436 15997
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 18788 16056 18840 16108
rect 9312 15852 9364 15904
rect 11428 15852 11480 15904
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 12992 15852 13044 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 14556 15852 14608 15904
rect 16028 15852 16080 15904
rect 16304 15895 16356 15904
rect 16304 15861 16313 15895
rect 16313 15861 16347 15895
rect 16347 15861 16356 15895
rect 16304 15852 16356 15861
rect 16396 15852 16448 15904
rect 16948 15852 17000 15904
rect 19616 15988 19668 16040
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 11888 15648 11940 15700
rect 16212 15648 16264 15700
rect 17224 15648 17276 15700
rect 17684 15648 17736 15700
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 10784 15580 10836 15632
rect 12624 15623 12676 15632
rect 8760 15512 8812 15564
rect 8944 15512 8996 15564
rect 11244 15512 11296 15564
rect 11336 15512 11388 15564
rect 12624 15589 12633 15623
rect 12633 15589 12667 15623
rect 12667 15589 12676 15623
rect 12624 15580 12676 15589
rect 15384 15623 15436 15632
rect 15384 15589 15393 15623
rect 15393 15589 15427 15623
rect 15427 15589 15436 15623
rect 15384 15580 15436 15589
rect 16580 15580 16632 15632
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 13544 15512 13596 15564
rect 16304 15512 16356 15564
rect 9036 15444 9088 15496
rect 9220 15444 9272 15496
rect 9956 15444 10008 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 10876 15308 10928 15360
rect 11980 15444 12032 15496
rect 13084 15444 13136 15496
rect 15384 15444 15436 15496
rect 15660 15444 15712 15496
rect 16764 15444 16816 15496
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 12808 15419 12860 15428
rect 12808 15385 12817 15419
rect 12817 15385 12851 15419
rect 12851 15385 12860 15419
rect 12808 15376 12860 15385
rect 17224 15376 17276 15428
rect 17960 15376 18012 15428
rect 13268 15308 13320 15360
rect 15200 15308 15252 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9956 15104 10008 15156
rect 10416 15147 10468 15156
rect 10416 15113 10425 15147
rect 10425 15113 10459 15147
rect 10459 15113 10468 15147
rect 10416 15104 10468 15113
rect 11888 15104 11940 15156
rect 12256 15104 12308 15156
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 9128 14968 9180 15020
rect 10324 15011 10376 15020
rect 10324 14977 10366 15011
rect 10366 14977 10376 15011
rect 10324 14968 10376 14977
rect 11704 14968 11756 15020
rect 11796 14968 11848 15020
rect 12532 14968 12584 15020
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 15108 15104 15160 15156
rect 15752 15104 15804 15156
rect 16580 15036 16632 15088
rect 13544 14968 13596 15020
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14464 15011 14516 15020
rect 14280 14968 14332 14977
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 16396 14968 16448 15020
rect 16488 14968 16540 15020
rect 17684 15011 17736 15020
rect 17684 14977 17693 15011
rect 17693 14977 17727 15011
rect 17727 14977 17736 15011
rect 17684 14968 17736 14977
rect 13728 14900 13780 14952
rect 10048 14832 10100 14884
rect 12624 14832 12676 14884
rect 15200 14943 15252 14952
rect 15200 14909 15209 14943
rect 15209 14909 15243 14943
rect 15243 14909 15252 14943
rect 15200 14900 15252 14909
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 15292 14832 15344 14884
rect 15844 14900 15896 14952
rect 17776 14900 17828 14952
rect 16764 14832 16816 14884
rect 18236 14832 18288 14884
rect 10232 14807 10284 14816
rect 10232 14773 10241 14807
rect 10241 14773 10275 14807
rect 10275 14773 10284 14807
rect 10232 14764 10284 14773
rect 12348 14807 12400 14816
rect 12348 14773 12357 14807
rect 12357 14773 12391 14807
rect 12391 14773 12400 14807
rect 12348 14764 12400 14773
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 13820 14764 13872 14816
rect 14004 14807 14056 14816
rect 14004 14773 14013 14807
rect 14013 14773 14047 14807
rect 14047 14773 14056 14807
rect 14004 14764 14056 14773
rect 15384 14764 15436 14816
rect 17776 14764 17828 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 9128 14603 9180 14612
rect 9128 14569 9137 14603
rect 9137 14569 9171 14603
rect 9171 14569 9180 14603
rect 9128 14560 9180 14569
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 12164 14560 12216 14612
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 12900 14560 12952 14612
rect 13912 14560 13964 14612
rect 14464 14603 14516 14612
rect 14464 14569 14473 14603
rect 14473 14569 14507 14603
rect 14507 14569 14516 14603
rect 14464 14560 14516 14569
rect 15568 14560 15620 14612
rect 17684 14560 17736 14612
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 1952 14424 2004 14476
rect 9312 14492 9364 14544
rect 10232 14424 10284 14476
rect 10324 14424 10376 14476
rect 14004 14492 14056 14544
rect 17316 14492 17368 14544
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 10508 14356 10560 14408
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 12808 14424 12860 14476
rect 13176 14424 13228 14476
rect 13544 14424 13596 14476
rect 18052 14467 18104 14476
rect 11796 14356 11848 14408
rect 13084 14356 13136 14408
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13728 14399 13780 14408
rect 13452 14356 13504 14365
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14372 14399 14424 14408
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 18052 14433 18061 14467
rect 18061 14433 18095 14467
rect 18095 14433 18104 14467
rect 18052 14424 18104 14433
rect 18236 14424 18288 14476
rect 16948 14356 17000 14365
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 20076 14356 20128 14408
rect 18604 14288 18656 14340
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 16488 14220 16540 14272
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9864 14016 9916 14068
rect 10416 14016 10468 14068
rect 15016 14016 15068 14068
rect 15568 14016 15620 14068
rect 10876 13948 10928 14000
rect 1952 13880 2004 13932
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 10968 13880 11020 13932
rect 11796 13880 11848 13932
rect 12808 13948 12860 14000
rect 17040 13948 17092 14000
rect 13176 13880 13228 13932
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 16948 13880 17000 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 17224 13880 17276 13932
rect 12348 13812 12400 13864
rect 12624 13787 12676 13796
rect 12624 13753 12633 13787
rect 12633 13753 12667 13787
rect 12667 13753 12676 13787
rect 12624 13744 12676 13753
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 9864 13676 9916 13728
rect 10784 13676 10836 13728
rect 11612 13676 11664 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10968 13472 11020 13524
rect 13544 13472 13596 13524
rect 14372 13472 14424 13524
rect 16948 13472 17000 13524
rect 8208 13336 8260 13388
rect 10508 13336 10560 13388
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 15016 13268 15068 13320
rect 15936 13311 15988 13320
rect 15936 13277 15970 13311
rect 15970 13277 15988 13311
rect 9956 13200 10008 13252
rect 14740 13243 14792 13252
rect 14740 13209 14749 13243
rect 14749 13209 14783 13243
rect 14783 13209 14792 13243
rect 14740 13200 14792 13209
rect 15200 13200 15252 13252
rect 15936 13268 15988 13277
rect 17132 13200 17184 13252
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 10876 12971 10928 12980
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 13452 12928 13504 12980
rect 14740 12928 14792 12980
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 18604 12971 18656 12980
rect 18604 12937 18613 12971
rect 18613 12937 18647 12971
rect 18647 12937 18656 12971
rect 18604 12928 18656 12937
rect 10600 12860 10652 12912
rect 15292 12903 15344 12912
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 10508 12792 10560 12844
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 13268 12792 13320 12844
rect 12808 12724 12860 12776
rect 13544 12792 13596 12844
rect 15292 12869 15301 12903
rect 15301 12869 15335 12903
rect 15335 12869 15344 12903
rect 15292 12860 15344 12869
rect 15016 12792 15068 12844
rect 15568 12835 15620 12844
rect 15568 12801 15577 12835
rect 15577 12801 15611 12835
rect 15611 12801 15620 12835
rect 15568 12792 15620 12801
rect 19340 12792 19392 12844
rect 38292 12835 38344 12844
rect 38292 12801 38301 12835
rect 38301 12801 38335 12835
rect 38335 12801 38344 12835
rect 38292 12792 38344 12801
rect 16488 12724 16540 12776
rect 13728 12656 13780 12708
rect 16580 12656 16632 12708
rect 17040 12656 17092 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 6552 12316 6604 12368
rect 17040 12291 17092 12300
rect 17040 12257 17049 12291
rect 17049 12257 17083 12291
rect 17083 12257 17092 12291
rect 17040 12248 17092 12257
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6944 1636 6996
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 37556 5695 37608 5704
rect 37556 5661 37565 5695
rect 37565 5661 37599 5695
rect 37599 5661 37608 5695
rect 37556 5652 37608 5661
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 9128 3068 9180 3120
rect 9036 2864 9088 2916
rect 37556 2864 37608 2916
rect 25872 2796 25924 2848
rect 32312 2839 32364 2848
rect 32312 2805 32321 2839
rect 32321 2805 32355 2839
rect 32355 2805 32364 2839
rect 32312 2796 32364 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 19340 2592 19392 2644
rect 15292 2456 15344 2508
rect 20 2388 72 2440
rect 6460 2388 6512 2440
rect 19432 2456 19484 2508
rect 24768 2456 24820 2508
rect 19340 2388 19392 2440
rect 25872 2431 25924 2440
rect 25872 2397 25881 2431
rect 25881 2397 25915 2431
rect 25915 2397 25924 2431
rect 25872 2388 25924 2397
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 12900 2252 12952 2304
rect 25780 2252 25832 2304
rect 32220 2252 32272 2304
rect 38660 2252 38712 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 39200 718 39800
rect 7102 39200 7158 39800
rect 13542 39200 13598 39800
rect 19982 39200 20038 39800
rect 26422 39200 26478 39800
rect 32862 39200 32918 39800
rect 39302 39200 39358 39800
rect 676 37262 704 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 7116 37330 7144 39200
rect 13556 37346 13584 39200
rect 7104 37324 7156 37330
rect 13556 37318 13676 37346
rect 7104 37266 7156 37272
rect 664 37256 716 37262
rect 664 37198 716 37204
rect 13648 37210 13676 37318
rect 19996 37262 20024 39200
rect 19432 37256 19484 37262
rect 7104 37188 7156 37194
rect 13648 37182 13860 37210
rect 19432 37198 19484 37204
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 7104 37130 7156 37136
rect 3792 37120 3844 37126
rect 3792 37062 3844 37068
rect 1676 34604 1728 34610
rect 1676 34546 1728 34552
rect 1688 28150 1716 34546
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34105 1808 34342
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2504 31748 2556 31754
rect 2504 31690 2556 31696
rect 2516 31278 2544 31690
rect 2792 31414 2820 31758
rect 2780 31408 2832 31414
rect 2780 31350 2832 31356
rect 3804 31346 3832 37062
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 6828 32428 6880 32434
rect 6828 32370 6880 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 6368 31952 6420 31958
rect 6368 31894 6420 31900
rect 6460 31952 6512 31958
rect 6460 31894 6512 31900
rect 5172 31816 5224 31822
rect 5172 31758 5224 31764
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 3792 31340 3844 31346
rect 3792 31282 3844 31288
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 1952 31272 2004 31278
rect 1952 31214 2004 31220
rect 2504 31272 2556 31278
rect 2504 31214 2556 31220
rect 2596 31272 2648 31278
rect 2596 31214 2648 31220
rect 1676 28144 1728 28150
rect 1676 28086 1728 28092
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1596 26382 1624 27950
rect 1860 27464 1912 27470
rect 1860 27406 1912 27412
rect 1768 27328 1820 27334
rect 1766 27296 1768 27305
rect 1820 27296 1822 27305
rect 1766 27231 1822 27240
rect 1872 27130 1900 27406
rect 1860 27124 1912 27130
rect 1860 27066 1912 27072
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 24750 1624 26318
rect 1584 24744 1636 24750
rect 1584 24686 1636 24692
rect 1596 24274 1624 24686
rect 1584 24268 1636 24274
rect 1584 24210 1636 24216
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 1780 20505 1808 20742
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19242 1900 19654
rect 1964 19446 1992 31214
rect 2608 30802 2636 31214
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 2596 30796 2648 30802
rect 2596 30738 2648 30744
rect 2136 30728 2188 30734
rect 2136 30670 2188 30676
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 2148 30190 2176 30670
rect 4436 30592 4488 30598
rect 4436 30534 4488 30540
rect 4448 30394 4476 30534
rect 4436 30388 4488 30394
rect 4436 30330 4488 30336
rect 4620 30320 4672 30326
rect 4620 30262 4672 30268
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 4068 30252 4120 30258
rect 4068 30194 4120 30200
rect 2136 30184 2188 30190
rect 2136 30126 2188 30132
rect 2148 28014 2176 30126
rect 2700 29850 2728 30194
rect 3884 30048 3936 30054
rect 3884 29990 3936 29996
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 3896 29714 3924 29990
rect 4080 29850 4108 30194
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29844 4120 29850
rect 4068 29786 4120 29792
rect 4160 29844 4212 29850
rect 4160 29786 4212 29792
rect 3884 29708 3936 29714
rect 3884 29650 3936 29656
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 2136 28008 2188 28014
rect 2136 27950 2188 27956
rect 2424 27674 2452 28018
rect 2412 27668 2464 27674
rect 2412 27610 2464 27616
rect 2700 27470 2728 29582
rect 3516 29164 3568 29170
rect 3516 29106 3568 29112
rect 3528 28218 3556 29106
rect 4172 29050 4200 29786
rect 4632 29714 4660 30262
rect 4620 29708 4672 29714
rect 4620 29650 4672 29656
rect 4816 29578 4844 30670
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4080 29034 4200 29050
rect 4896 29096 4948 29102
rect 5000 29050 5028 31282
rect 5184 30054 5212 31758
rect 5448 31748 5500 31754
rect 5368 31708 5448 31736
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 5368 29646 5396 31708
rect 5448 31690 5500 31696
rect 5828 31482 5856 31758
rect 5908 31680 5960 31686
rect 5908 31622 5960 31628
rect 6000 31680 6052 31686
rect 6000 31622 6052 31628
rect 5816 31476 5868 31482
rect 5816 31418 5868 31424
rect 5724 31136 5776 31142
rect 5724 31078 5776 31084
rect 5736 30802 5764 31078
rect 5724 30796 5776 30802
rect 5724 30738 5776 30744
rect 5448 30728 5500 30734
rect 5448 30670 5500 30676
rect 5460 29714 5488 30670
rect 5448 29708 5500 29714
rect 5448 29650 5500 29656
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5368 29102 5396 29582
rect 4948 29044 5028 29050
rect 4896 29038 5028 29044
rect 5356 29096 5408 29102
rect 5356 29038 5408 29044
rect 4080 29028 4212 29034
rect 4080 29022 4160 29028
rect 4080 28642 4108 29022
rect 4908 29022 5028 29038
rect 4160 28970 4212 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4896 28756 4948 28762
rect 4896 28698 4948 28704
rect 4080 28614 4200 28642
rect 4172 28558 4200 28614
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 3976 28416 4028 28422
rect 3976 28358 4028 28364
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 3988 28082 4016 28358
rect 3976 28076 4028 28082
rect 3976 28018 4028 28024
rect 4172 27962 4200 28494
rect 4620 28212 4672 28218
rect 4620 28154 4672 28160
rect 4080 27934 4200 27962
rect 4080 27656 4108 27934
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4080 27628 4200 27656
rect 2688 27464 2740 27470
rect 2688 27406 2740 27412
rect 2042 27024 2098 27033
rect 2042 26959 2044 26968
rect 2096 26959 2098 26968
rect 2044 26930 2096 26936
rect 2596 26308 2648 26314
rect 2596 26250 2648 26256
rect 2608 26042 2636 26250
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 2700 25906 2728 27406
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 3332 26784 3384 26790
rect 3332 26726 3384 26732
rect 3344 25974 3372 26726
rect 3528 26518 3556 26930
rect 3516 26512 3568 26518
rect 3516 26454 3568 26460
rect 3620 26314 3648 26930
rect 3884 26920 3936 26926
rect 3884 26862 3936 26868
rect 3896 26382 3924 26862
rect 3988 26586 4016 27338
rect 4172 26874 4200 27628
rect 4632 27606 4660 28154
rect 4804 28008 4856 28014
rect 4804 27950 4856 27956
rect 4712 27940 4764 27946
rect 4712 27882 4764 27888
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4632 27470 4660 27542
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4724 27062 4752 27882
rect 4816 27674 4844 27950
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4908 27538 4936 28698
rect 4896 27532 4948 27538
rect 4896 27474 4948 27480
rect 5000 27402 5028 29022
rect 5264 28756 5316 28762
rect 5264 28698 5316 28704
rect 5276 28506 5304 28698
rect 5368 28558 5396 29038
rect 5092 28478 5304 28506
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5092 27470 5120 28478
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5172 28008 5224 28014
rect 5172 27950 5224 27956
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 4988 27396 5040 27402
rect 4988 27338 5040 27344
rect 4712 27056 4764 27062
rect 4712 26998 4764 27004
rect 4080 26846 4200 26874
rect 3976 26580 4028 26586
rect 3976 26522 4028 26528
rect 4080 26466 4108 26846
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26466 4660 26726
rect 4080 26438 4200 26466
rect 4172 26382 4200 26438
rect 4540 26438 4660 26466
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 4160 26376 4212 26382
rect 4160 26318 4212 26324
rect 3608 26308 3660 26314
rect 3608 26250 3660 26256
rect 4436 26308 4488 26314
rect 4436 26250 4488 26256
rect 3332 25968 3384 25974
rect 3332 25910 3384 25916
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 2700 24818 2728 25842
rect 4080 25498 4108 25842
rect 4448 25786 4476 26250
rect 4540 25974 4568 26438
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 4632 26042 4660 26318
rect 4620 26036 4672 26042
rect 4620 25978 4672 25984
rect 4528 25968 4580 25974
rect 4528 25910 4580 25916
rect 4448 25758 4660 25786
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 3148 24812 3200 24818
rect 3148 24754 3200 24760
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 2240 24206 2268 24550
rect 2332 24410 2360 24754
rect 2320 24404 2372 24410
rect 2320 24346 2372 24352
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2424 23712 2452 24754
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 2332 23684 2452 23712
rect 2332 22234 2360 23684
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2688 22500 2740 22506
rect 2688 22442 2740 22448
rect 2320 22228 2372 22234
rect 2320 22170 2372 22176
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 2148 21622 2176 21966
rect 2136 21616 2188 21622
rect 2136 21558 2188 21564
rect 2332 20466 2360 22170
rect 2700 22030 2728 22442
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2792 21690 2820 22578
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2884 21554 2912 22374
rect 2976 22030 3004 22578
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 2872 21548 2924 21554
rect 2872 21490 2924 21496
rect 3068 21486 3096 24550
rect 3160 24206 3188 24754
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3424 24336 3476 24342
rect 3424 24278 3476 24284
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3252 23730 3280 23802
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3436 23662 3464 24278
rect 3620 23798 3648 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24290 4660 25758
rect 4724 25294 4752 26998
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 4804 26852 4856 26858
rect 4804 26794 4856 26800
rect 4816 26042 4844 26794
rect 4896 26784 4948 26790
rect 4896 26726 4948 26732
rect 4804 26036 4856 26042
rect 4804 25978 4856 25984
rect 4816 25294 4844 25978
rect 4908 25702 4936 26726
rect 5000 25770 5028 26930
rect 5092 26518 5120 27406
rect 5184 27062 5212 27950
rect 5276 27946 5304 28358
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 5172 27056 5224 27062
rect 5172 26998 5224 27004
rect 5276 26994 5304 27882
rect 5368 27130 5396 28154
rect 5460 27878 5488 29650
rect 5540 29640 5592 29646
rect 5540 29582 5592 29588
rect 5552 28218 5580 29582
rect 5540 28212 5592 28218
rect 5540 28154 5592 28160
rect 5736 28082 5764 30738
rect 5816 30592 5868 30598
rect 5816 30534 5868 30540
rect 5828 30394 5856 30534
rect 5816 30388 5868 30394
rect 5816 30330 5868 30336
rect 5816 30048 5868 30054
rect 5816 29990 5868 29996
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5644 27606 5672 28018
rect 5632 27600 5684 27606
rect 5632 27542 5684 27548
rect 5448 27396 5500 27402
rect 5448 27338 5500 27344
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 5368 26994 5396 27066
rect 5264 26988 5316 26994
rect 5264 26930 5316 26936
rect 5356 26988 5408 26994
rect 5356 26930 5408 26936
rect 5080 26512 5132 26518
rect 5080 26454 5132 26460
rect 5092 26382 5120 26454
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 4988 25764 5040 25770
rect 4988 25706 5040 25712
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 5184 24698 5212 26386
rect 5276 25974 5304 26930
rect 5368 26246 5396 26930
rect 5460 26586 5488 27338
rect 5540 27056 5592 27062
rect 5540 26998 5592 27004
rect 5448 26580 5500 26586
rect 5448 26522 5500 26528
rect 5552 26518 5580 26998
rect 5828 26994 5856 29990
rect 5920 29714 5948 31622
rect 6012 31346 6040 31622
rect 6000 31340 6052 31346
rect 6000 31282 6052 31288
rect 6380 30258 6408 31894
rect 6472 31822 6500 31894
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6472 31278 6500 31758
rect 6656 31346 6684 31758
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6644 31340 6696 31346
rect 6644 31282 6696 31288
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 6552 31204 6604 31210
rect 6552 31146 6604 31152
rect 6564 30394 6592 31146
rect 6644 30864 6696 30870
rect 6644 30806 6696 30812
rect 6552 30388 6604 30394
rect 6552 30330 6604 30336
rect 6656 30258 6684 30806
rect 6748 30802 6776 31418
rect 6736 30796 6788 30802
rect 6736 30738 6788 30744
rect 6840 30326 6868 32370
rect 6828 30320 6880 30326
rect 6828 30262 6880 30268
rect 6368 30252 6420 30258
rect 6368 30194 6420 30200
rect 6644 30252 6696 30258
rect 6644 30194 6696 30200
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 6656 28370 6684 29990
rect 6748 29170 6776 30126
rect 6840 30054 6868 30126
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6828 29572 6880 29578
rect 6828 29514 6880 29520
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 6736 29164 6788 29170
rect 6736 29106 6788 29112
rect 6748 28490 6776 29106
rect 6840 28558 6868 29514
rect 7024 29306 7052 29514
rect 7012 29300 7064 29306
rect 7012 29242 7064 29248
rect 7024 28994 7052 29242
rect 6932 28966 7052 28994
rect 6932 28694 6960 28966
rect 6920 28688 6972 28694
rect 6920 28630 6972 28636
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6736 28484 6788 28490
rect 6736 28426 6788 28432
rect 6656 28342 6868 28370
rect 6092 28144 6144 28150
rect 6092 28086 6144 28092
rect 5816 26988 5868 26994
rect 5816 26930 5868 26936
rect 5540 26512 5592 26518
rect 5540 26454 5592 26460
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 5368 25838 5396 26182
rect 5552 25906 5580 26454
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5356 25832 5408 25838
rect 5356 25774 5408 25780
rect 5368 25226 5396 25774
rect 5736 25770 5764 26250
rect 5724 25764 5776 25770
rect 5724 25706 5776 25712
rect 5632 25424 5684 25430
rect 5736 25412 5764 25706
rect 5684 25384 5764 25412
rect 5632 25366 5684 25372
rect 5356 25220 5408 25226
rect 5356 25162 5408 25168
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5276 24886 5304 25094
rect 5264 24880 5316 24886
rect 5264 24822 5316 24828
rect 5184 24670 5304 24698
rect 5276 24614 5304 24670
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 4540 24262 4660 24290
rect 4908 24274 4936 24550
rect 4896 24268 4948 24274
rect 4436 24200 4488 24206
rect 4436 24142 4488 24148
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 3608 23792 3660 23798
rect 3608 23734 3660 23740
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3436 23066 3464 23598
rect 3436 23038 3556 23066
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3436 22710 3464 22918
rect 3424 22704 3476 22710
rect 3424 22646 3476 22652
rect 3332 22432 3384 22438
rect 3332 22374 3384 22380
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2320 20460 2372 20466
rect 2320 20402 2372 20408
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 2148 19854 2176 20198
rect 2240 20058 2268 20402
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2976 19990 3004 20810
rect 3068 20534 3096 21422
rect 3252 20942 3280 21830
rect 3344 21486 3372 22374
rect 3436 22030 3464 22646
rect 3528 22642 3556 23038
rect 3712 22778 3740 23802
rect 4448 23526 4476 24142
rect 4540 24070 4568 24262
rect 4896 24210 4948 24216
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4632 23662 4660 24142
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4724 23186 4752 23666
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4816 23254 4844 23462
rect 4804 23248 4856 23254
rect 4804 23190 4856 23196
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3528 22166 3556 22578
rect 3516 22160 3568 22166
rect 3516 22102 3568 22108
rect 3712 22094 3740 22714
rect 4356 22642 4384 23122
rect 4908 23066 4936 24210
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 4724 23038 4936 23066
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4160 22500 4212 22506
rect 4080 22460 4160 22488
rect 4080 22098 4108 22460
rect 4160 22442 4212 22448
rect 4356 22438 4384 22578
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3620 22066 3740 22094
rect 4068 22092 4120 22098
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3620 21962 3648 22066
rect 4068 22034 4120 22040
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 4264 21690 4292 21966
rect 4252 21684 4304 21690
rect 4252 21626 4304 21632
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3056 20528 3108 20534
rect 3056 20470 3108 20476
rect 3436 20398 3464 20742
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3056 20324 3108 20330
rect 3056 20266 3108 20272
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 1952 19440 2004 19446
rect 1952 19382 2004 19388
rect 2976 19310 3004 19926
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 1860 19236 1912 19242
rect 1860 19178 1912 19184
rect 1872 17134 1900 19178
rect 2976 18766 3004 19246
rect 3068 18834 3096 20266
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3252 19922 3280 20198
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 3068 18222 3096 18770
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3160 17610 3188 19314
rect 3252 18970 3280 19858
rect 3436 19854 3464 20334
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3896 18154 3924 20402
rect 3988 20398 4016 20878
rect 4264 20466 4292 20946
rect 4632 20618 4660 22578
rect 4724 21554 4752 23038
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4816 21486 4844 22578
rect 4908 22166 4936 22918
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 4896 22160 4948 22166
rect 4896 22102 4948 22108
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4632 20590 4752 20618
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 3988 19514 4016 20334
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 19718 4108 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4632 19174 4660 20402
rect 4724 19530 4752 20590
rect 4816 20058 4844 21422
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4908 19786 4936 21966
rect 5000 21622 5028 22510
rect 4988 21616 5040 21622
rect 4988 21558 5040 21564
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4724 19502 4844 19530
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4448 18290 4476 18702
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4632 18290 4660 18566
rect 4724 18426 4752 19382
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4448 18170 4476 18226
rect 4816 18170 4844 19502
rect 3884 18148 3936 18154
rect 4448 18142 4660 18170
rect 3884 18090 3936 18096
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18142
rect 4724 18142 4844 18170
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4724 17678 4752 18142
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4816 17678 4844 18022
rect 5184 17678 5212 23122
rect 5368 23118 5396 24006
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5448 22568 5500 22574
rect 5736 22556 5764 25384
rect 5828 22710 5856 26930
rect 5908 26784 5960 26790
rect 5908 26726 5960 26732
rect 5920 26450 5948 26726
rect 5908 26444 5960 26450
rect 5908 26386 5960 26392
rect 6104 25430 6132 28086
rect 6460 27056 6512 27062
rect 6460 26998 6512 27004
rect 6184 26988 6236 26994
rect 6184 26930 6236 26936
rect 6196 26586 6224 26930
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6472 26382 6500 26998
rect 6840 26382 6868 28342
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6460 25900 6512 25906
rect 6460 25842 6512 25848
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 5908 25424 5960 25430
rect 5908 25366 5960 25372
rect 6092 25424 6144 25430
rect 6092 25366 6144 25372
rect 5920 22778 5948 25366
rect 6472 25226 6500 25842
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6092 25152 6144 25158
rect 6092 25094 6144 25100
rect 6000 24676 6052 24682
rect 6000 24618 6052 24624
rect 6012 24274 6040 24618
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 6104 24206 6132 25094
rect 6472 24818 6500 25162
rect 6656 25158 6684 25774
rect 6748 25498 6776 25842
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6460 24812 6512 24818
rect 6460 24754 6512 24760
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 6012 23866 6040 24074
rect 6104 23866 6132 24142
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 5816 22704 5868 22710
rect 5816 22646 5868 22652
rect 5736 22528 5856 22556
rect 5448 22510 5500 22516
rect 5460 22030 5488 22510
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5644 21554 5672 21898
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5644 21026 5672 21490
rect 5552 20998 5672 21026
rect 5552 20618 5580 20998
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5460 20590 5580 20618
rect 5460 20534 5488 20590
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5276 19378 5304 20402
rect 5460 19514 5488 20470
rect 5644 20262 5672 20878
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5276 17678 5304 19314
rect 5460 19310 5488 19450
rect 5644 19378 5672 20198
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5552 18766 5580 19178
rect 5644 18970 5672 19314
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5552 17746 5580 18226
rect 5736 18222 5764 19722
rect 5828 18680 5856 22528
rect 6104 22166 6132 23054
rect 6472 22642 6500 24754
rect 6748 24138 6776 25434
rect 6840 25294 6868 26318
rect 7116 25906 7144 37130
rect 13832 37126 13860 37182
rect 13820 37120 13872 37126
rect 13820 37062 13872 37068
rect 19444 36922 19472 37198
rect 26436 37126 26464 39200
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 20076 37120 20128 37126
rect 20076 37062 20128 37068
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 20088 36786 20116 37062
rect 20076 36780 20128 36786
rect 20076 36722 20128 36728
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 17316 34128 17368 34134
rect 17316 34070 17368 34076
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 12624 33992 12676 33998
rect 12624 33934 12676 33940
rect 9680 33856 9732 33862
rect 9680 33798 9732 33804
rect 9692 33590 9720 33798
rect 9680 33584 9732 33590
rect 9680 33526 9732 33532
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 8116 33312 8168 33318
rect 8116 33254 8168 33260
rect 7472 32904 7524 32910
rect 7472 32846 7524 32852
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 7300 31346 7328 32506
rect 7288 31340 7340 31346
rect 7288 31282 7340 31288
rect 7300 29646 7328 31282
rect 7380 30660 7432 30666
rect 7380 30602 7432 30608
rect 7288 29640 7340 29646
rect 7288 29582 7340 29588
rect 7196 29504 7248 29510
rect 7196 29446 7248 29452
rect 7208 28626 7236 29446
rect 7196 28620 7248 28626
rect 7196 28562 7248 28568
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7300 26314 7328 28494
rect 7288 26308 7340 26314
rect 7288 26250 7340 26256
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 7024 24410 7052 25638
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6552 23248 6604 23254
rect 6552 23190 6604 23196
rect 6564 22710 6592 23190
rect 6552 22704 6604 22710
rect 6552 22646 6604 22652
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6092 22160 6144 22166
rect 6092 22102 6144 22108
rect 6104 21486 6132 22102
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 21554 6684 21830
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 6012 20942 6040 21354
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6276 21072 6328 21078
rect 6748 21049 6776 21082
rect 7024 21078 7052 24210
rect 7116 24206 7144 25094
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7116 21146 7144 23054
rect 7208 22094 7236 25230
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7300 24070 7328 25094
rect 7288 24064 7340 24070
rect 7288 24006 7340 24012
rect 7300 23730 7328 24006
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7208 22066 7328 22094
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7012 21072 7064 21078
rect 6276 21014 6328 21020
rect 6734 21040 6790 21049
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 5920 20602 5948 20878
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 6104 20466 6132 20810
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 5908 18692 5960 18698
rect 5828 18652 5908 18680
rect 5908 18634 5960 18640
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 3148 17604 3200 17610
rect 3148 17546 3200 17552
rect 5184 17270 5212 17614
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 4080 16794 4108 17138
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 5368 16590 5396 17478
rect 5552 17338 5580 17682
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 6012 16590 6040 19382
rect 6104 18358 6132 20266
rect 6288 20058 6316 21014
rect 7012 21014 7064 21020
rect 6734 20975 6790 20984
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6288 18426 6316 19994
rect 6380 19854 6408 20878
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6472 19922 6500 20538
rect 6564 20058 6592 20878
rect 6932 20618 6960 20878
rect 7024 20806 7052 21014
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 6840 20590 6960 20618
rect 6840 20398 6868 20590
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6564 19378 6592 19790
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6656 18834 6684 19314
rect 7300 19310 7328 22066
rect 7392 21690 7420 30602
rect 7484 28762 7512 32846
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7668 32434 7696 32710
rect 8128 32502 8156 33254
rect 8312 32570 8340 33458
rect 8852 33312 8904 33318
rect 8852 33254 8904 33260
rect 8864 32978 8892 33254
rect 9876 33114 9904 33934
rect 12636 33522 12664 33934
rect 12900 33924 12952 33930
rect 12900 33866 12952 33872
rect 12624 33516 12676 33522
rect 12624 33458 12676 33464
rect 12072 33448 12124 33454
rect 12072 33390 12124 33396
rect 10968 33312 11020 33318
rect 10968 33254 11020 33260
rect 9864 33108 9916 33114
rect 9864 33050 9916 33056
rect 8852 32972 8904 32978
rect 8852 32914 8904 32920
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8300 32564 8352 32570
rect 8300 32506 8352 32512
rect 8116 32496 8168 32502
rect 8116 32438 8168 32444
rect 7656 32428 7708 32434
rect 7656 32370 7708 32376
rect 7932 32224 7984 32230
rect 7932 32166 7984 32172
rect 7944 31958 7972 32166
rect 7932 31952 7984 31958
rect 7932 31894 7984 31900
rect 7748 31136 7800 31142
rect 7748 31078 7800 31084
rect 7760 30734 7788 31078
rect 7748 30728 7800 30734
rect 7748 30670 7800 30676
rect 7564 30320 7616 30326
rect 7564 30262 7616 30268
rect 7576 30122 7604 30262
rect 7564 30116 7616 30122
rect 7564 30058 7616 30064
rect 7944 30054 7972 31894
rect 8024 31816 8076 31822
rect 8024 31758 8076 31764
rect 8036 31346 8064 31758
rect 8128 31482 8156 32438
rect 8300 31748 8352 31754
rect 8300 31690 8352 31696
rect 8116 31476 8168 31482
rect 8116 31418 8168 31424
rect 8024 31340 8076 31346
rect 8024 31282 8076 31288
rect 8024 31136 8076 31142
rect 8024 31078 8076 31084
rect 8036 30734 8064 31078
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 8036 29850 8064 30126
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 8128 29714 8156 31418
rect 8312 31346 8340 31690
rect 8297 31340 8349 31346
rect 8297 31282 8349 31288
rect 8312 30802 8340 31282
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8116 29708 8168 29714
rect 8116 29650 8168 29656
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 7472 28756 7524 28762
rect 7472 28698 7524 28704
rect 8024 28552 8076 28558
rect 8024 28494 8076 28500
rect 8036 28218 8064 28494
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 8024 28212 8076 28218
rect 8024 28154 8076 28160
rect 7656 28144 7708 28150
rect 7656 28086 7708 28092
rect 7668 26058 7696 28086
rect 7852 27674 7880 28154
rect 8220 28014 8248 29582
rect 8404 29306 8432 32846
rect 8760 32564 8812 32570
rect 8760 32506 8812 32512
rect 8576 32292 8628 32298
rect 8576 32234 8628 32240
rect 8588 31958 8616 32234
rect 8668 32020 8720 32026
rect 8668 31962 8720 31968
rect 8576 31952 8628 31958
rect 8576 31894 8628 31900
rect 8680 31346 8708 31962
rect 8668 31340 8720 31346
rect 8668 31282 8720 31288
rect 8576 31204 8628 31210
rect 8576 31146 8628 31152
rect 8484 30796 8536 30802
rect 8484 30738 8536 30744
rect 8496 30394 8524 30738
rect 8588 30598 8616 31146
rect 8576 30592 8628 30598
rect 8576 30534 8628 30540
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 8680 29594 8708 31282
rect 8772 31278 8800 32506
rect 8864 32366 8892 32914
rect 10980 32910 11008 33254
rect 9404 32904 9456 32910
rect 9404 32846 9456 32852
rect 10968 32904 11020 32910
rect 10968 32846 11020 32852
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 8852 32360 8904 32366
rect 8852 32302 8904 32308
rect 9416 32026 9444 32846
rect 10324 32768 10376 32774
rect 10324 32710 10376 32716
rect 10336 32502 10364 32710
rect 10324 32496 10376 32502
rect 10324 32438 10376 32444
rect 9496 32428 9548 32434
rect 9496 32370 9548 32376
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9220 31952 9272 31958
rect 9220 31894 9272 31900
rect 8760 31272 8812 31278
rect 8760 31214 8812 31220
rect 9232 30258 9260 31894
rect 9508 31754 9536 32370
rect 10980 32366 11008 32846
rect 11072 32570 11100 32846
rect 11060 32564 11112 32570
rect 11060 32506 11112 32512
rect 11072 32434 11100 32506
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 10968 32360 11020 32366
rect 10968 32302 11020 32308
rect 9772 32292 9824 32298
rect 9772 32234 9824 32240
rect 11888 32292 11940 32298
rect 11888 32234 11940 32240
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 9416 31726 9536 31754
rect 9416 30326 9444 31726
rect 9496 31272 9548 31278
rect 9496 31214 9548 31220
rect 9508 30802 9536 31214
rect 9496 30796 9548 30802
rect 9496 30738 9548 30744
rect 9600 30734 9628 31758
rect 9692 31346 9720 31826
rect 9784 31414 9812 32234
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 9956 31680 10008 31686
rect 9956 31622 10008 31628
rect 9772 31408 9824 31414
rect 9772 31350 9824 31356
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9784 30598 9812 31350
rect 9864 31340 9916 31346
rect 9968 31328 9996 31622
rect 9916 31300 9996 31328
rect 9864 31282 9916 31288
rect 9862 30832 9918 30841
rect 9968 30802 9996 31300
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 10060 30870 10088 31078
rect 10048 30864 10100 30870
rect 10048 30806 10100 30812
rect 9862 30767 9918 30776
rect 9956 30796 10008 30802
rect 9876 30666 9904 30767
rect 9956 30738 10008 30744
rect 9864 30660 9916 30666
rect 9864 30602 9916 30608
rect 9772 30592 9824 30598
rect 9772 30534 9824 30540
rect 9968 30394 9996 30738
rect 10152 30734 10180 31758
rect 10336 30734 10364 31826
rect 10612 31822 10640 32166
rect 10980 31890 11008 32166
rect 11900 31890 11928 32234
rect 11980 32224 12032 32230
rect 11980 32166 12032 32172
rect 10968 31884 11020 31890
rect 11888 31884 11940 31890
rect 10968 31826 11020 31832
rect 11808 31844 11888 31872
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10692 31680 10744 31686
rect 10692 31622 10744 31628
rect 10704 31362 10732 31622
rect 10980 31414 11008 31826
rect 11060 31816 11112 31822
rect 11060 31758 11112 31764
rect 11152 31816 11204 31822
rect 11152 31758 11204 31764
rect 10784 31408 10836 31414
rect 10704 31356 10784 31362
rect 10704 31350 10836 31356
rect 10968 31408 11020 31414
rect 10968 31350 11020 31356
rect 10600 31340 10652 31346
rect 10600 31282 10652 31288
rect 10704 31334 10824 31350
rect 10612 30802 10640 31282
rect 10600 30796 10652 30802
rect 10600 30738 10652 30744
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10324 30728 10376 30734
rect 10324 30670 10376 30676
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 9956 30388 10008 30394
rect 9956 30330 10008 30336
rect 9404 30320 9456 30326
rect 9404 30262 9456 30268
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 9232 29782 9260 30194
rect 10612 30190 10640 30534
rect 10704 30394 10732 31334
rect 11072 30598 11100 31758
rect 11164 31278 11192 31758
rect 11244 31748 11296 31754
rect 11244 31690 11296 31696
rect 11256 31414 11284 31690
rect 11336 31680 11388 31686
rect 11336 31622 11388 31628
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11244 31408 11296 31414
rect 11244 31350 11296 31356
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 11244 31272 11296 31278
rect 11244 31214 11296 31220
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10692 30388 10744 30394
rect 10692 30330 10744 30336
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 9220 29776 9272 29782
rect 9220 29718 9272 29724
rect 10324 29708 10376 29714
rect 10324 29650 10376 29656
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 8496 29566 8708 29594
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 8760 29572 8812 29578
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 8312 28966 8340 29106
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 8404 28762 8432 29106
rect 8496 29034 8524 29566
rect 8760 29514 8812 29520
rect 8576 29504 8628 29510
rect 8576 29446 8628 29452
rect 8588 29238 8616 29446
rect 8576 29232 8628 29238
rect 8576 29174 8628 29180
rect 8668 29096 8720 29102
rect 8668 29038 8720 29044
rect 8484 29028 8536 29034
rect 8484 28970 8536 28976
rect 8392 28756 8444 28762
rect 8392 28698 8444 28704
rect 8496 28558 8524 28970
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 8496 27878 8524 28494
rect 8680 28218 8708 29038
rect 8772 28762 8800 29514
rect 9140 29102 9168 29582
rect 9324 29238 9352 29582
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9508 29238 9536 29446
rect 9312 29232 9364 29238
rect 9312 29174 9364 29180
rect 9496 29232 9548 29238
rect 9496 29174 9548 29180
rect 9128 29096 9180 29102
rect 9128 29038 9180 29044
rect 9496 29096 9548 29102
rect 9496 29038 9548 29044
rect 8760 28756 8812 28762
rect 8760 28698 8812 28704
rect 9404 28756 9456 28762
rect 9404 28698 9456 28704
rect 8772 28490 8800 28698
rect 8760 28484 8812 28490
rect 8760 28426 8812 28432
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 9416 28014 9444 28698
rect 9508 28218 9536 29038
rect 9600 28966 9628 29582
rect 10336 29170 10364 29650
rect 10324 29164 10376 29170
rect 10324 29106 10376 29112
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9600 28762 9628 28902
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 10520 28626 10548 29650
rect 10980 29646 11008 29990
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10600 29096 10652 29102
rect 10600 29038 10652 29044
rect 10508 28620 10560 28626
rect 10508 28562 10560 28568
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 7840 27668 7892 27674
rect 7840 27610 7892 27616
rect 8300 27600 8352 27606
rect 8300 27542 8352 27548
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7852 27130 7880 27406
rect 8208 27396 8260 27402
rect 8208 27338 8260 27344
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 8220 26994 8248 27338
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 7748 26852 7800 26858
rect 7748 26794 7800 26800
rect 7760 26450 7788 26794
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 8024 26240 8076 26246
rect 8024 26182 8076 26188
rect 7668 26030 7788 26058
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7392 20466 7420 21422
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7392 20058 7420 20402
rect 7484 20398 7512 25842
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7576 25294 7604 25638
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7484 19854 7512 20334
rect 7668 19922 7696 25842
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7760 19786 7788 26030
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 7944 24410 7972 24754
rect 8036 24750 8064 26182
rect 8312 25702 8340 27542
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8404 26314 8432 27270
rect 8588 26450 8616 27406
rect 9220 27396 9272 27402
rect 9220 27338 9272 27344
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 8668 26920 8720 26926
rect 8668 26862 8720 26868
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 8404 25498 8432 26250
rect 8588 26024 8616 26386
rect 8496 25996 8616 26024
rect 8392 25492 8444 25498
rect 8392 25434 8444 25440
rect 8496 25226 8524 25996
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8588 25498 8616 25842
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 8680 25294 8708 26862
rect 9232 26586 9260 27338
rect 9324 27130 9352 27338
rect 9312 27124 9364 27130
rect 9312 27066 9364 27072
rect 9416 26994 9444 27950
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9692 26926 9720 28494
rect 10520 28150 10548 28562
rect 10612 28558 10640 29038
rect 10704 28558 10732 29446
rect 10796 29306 10824 29582
rect 10784 29300 10836 29306
rect 10784 29242 10836 29248
rect 10966 29064 11022 29073
rect 10966 28999 10968 29008
rect 11020 28999 11022 29008
rect 10968 28970 11020 28976
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 9864 28144 9916 28150
rect 9864 28086 9916 28092
rect 10508 28144 10560 28150
rect 10508 28086 10560 28092
rect 9876 27402 9904 28086
rect 10980 28082 11008 28970
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 9864 27396 9916 27402
rect 9864 27338 9916 27344
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 8852 25900 8904 25906
rect 8852 25842 8904 25848
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 8484 25220 8536 25226
rect 8484 25162 8536 25168
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 8036 24274 8064 24686
rect 8772 24342 8800 25774
rect 8760 24336 8812 24342
rect 8760 24278 8812 24284
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 8036 23662 8064 24210
rect 8864 24138 8892 25842
rect 9232 25294 9260 26522
rect 9600 26382 9628 26862
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9692 26246 9720 26862
rect 9876 26353 9904 27338
rect 9862 26344 9918 26353
rect 9772 26308 9824 26314
rect 9862 26279 9918 26288
rect 9772 26250 9824 26256
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9692 25498 9720 25842
rect 9784 25770 9812 26250
rect 9876 26042 9904 26279
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9772 25764 9824 25770
rect 9772 25706 9824 25712
rect 9864 25764 9916 25770
rect 9864 25706 9916 25712
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9876 25430 9904 25706
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 9864 25424 9916 25430
rect 9864 25366 9916 25372
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9968 24818 9996 25230
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 9772 24676 9824 24682
rect 9772 24618 9824 24624
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 8116 24064 8168 24070
rect 8116 24006 8168 24012
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8128 23866 8156 24006
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8220 23798 8248 24006
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 8680 23322 8708 23666
rect 8864 23322 8892 24074
rect 9692 23798 9720 24550
rect 9784 23866 9812 24618
rect 9968 24206 9996 24754
rect 10060 24750 10088 25638
rect 10140 25152 10192 25158
rect 10428 25129 10456 28018
rect 10508 27668 10560 27674
rect 10508 27610 10560 27616
rect 10520 27334 10548 27610
rect 11164 27538 11192 31214
rect 11256 30784 11284 31214
rect 11348 31142 11376 31622
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11428 30796 11480 30802
rect 11256 30756 11428 30784
rect 11256 29850 11284 30756
rect 11428 30738 11480 30744
rect 11532 30734 11560 31622
rect 11704 30932 11756 30938
rect 11704 30874 11756 30880
rect 11612 30796 11664 30802
rect 11612 30738 11664 30744
rect 11520 30728 11572 30734
rect 11520 30670 11572 30676
rect 11532 30326 11560 30670
rect 11520 30320 11572 30326
rect 11520 30262 11572 30268
rect 11624 30258 11652 30738
rect 11612 30252 11664 30258
rect 11612 30194 11664 30200
rect 11244 29844 11296 29850
rect 11244 29786 11296 29792
rect 11716 29170 11744 30874
rect 11808 30734 11836 31844
rect 11888 31826 11940 31832
rect 11992 31754 12020 32166
rect 12084 31754 12112 33390
rect 12808 33312 12860 33318
rect 12808 33254 12860 33260
rect 12820 33114 12848 33254
rect 12912 33114 12940 33866
rect 13820 33516 13872 33522
rect 13820 33458 13872 33464
rect 12808 33108 12860 33114
rect 12808 33050 12860 33056
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 12912 32910 12940 33050
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 12716 32836 12768 32842
rect 12716 32778 12768 32784
rect 12728 32570 12756 32778
rect 12716 32564 12768 32570
rect 12716 32506 12768 32512
rect 12716 32428 12768 32434
rect 12716 32370 12768 32376
rect 12728 31890 12756 32370
rect 12716 31884 12768 31890
rect 12716 31826 12768 31832
rect 11980 31748 12032 31754
rect 12084 31726 12204 31754
rect 11980 31690 12032 31696
rect 12176 31414 12204 31726
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 12452 31482 12480 31622
rect 12440 31476 12492 31482
rect 12440 31418 12492 31424
rect 12164 31408 12216 31414
rect 12164 31350 12216 31356
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11900 30938 11928 31282
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12084 29714 12112 29786
rect 12072 29708 12124 29714
rect 12072 29650 12124 29656
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 11900 29170 11928 29514
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11152 27532 11204 27538
rect 11152 27474 11204 27480
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 10508 27328 10560 27334
rect 10508 27270 10560 27276
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 10520 25974 10548 27270
rect 11348 27062 11376 27270
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 10508 25968 10560 25974
rect 10508 25910 10560 25916
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10140 25094 10192 25100
rect 10414 25120 10470 25129
rect 10152 24886 10180 25094
rect 10414 25055 10470 25064
rect 10140 24880 10192 24886
rect 10140 24822 10192 24828
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9680 23792 9732 23798
rect 9680 23734 9732 23740
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8852 23316 8904 23322
rect 8852 23258 8904 23264
rect 8864 23118 8892 23258
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 8392 23044 8444 23050
rect 8392 22986 8444 22992
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7852 22438 7880 22918
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7852 22166 7880 22374
rect 7840 22160 7892 22166
rect 7840 22102 7892 22108
rect 8300 22160 8352 22166
rect 8300 22102 8352 22108
rect 7852 21554 7880 22102
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7852 21010 7880 21490
rect 7932 21412 7984 21418
rect 7932 21354 7984 21360
rect 7944 21146 7972 21354
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 8312 21078 8340 22102
rect 8404 21554 8432 22986
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8956 21554 8984 22034
rect 9416 21962 9444 22918
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9508 22094 9536 22578
rect 9600 22234 9628 23054
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 10060 22094 10088 24686
rect 10244 24410 10272 24754
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10232 23044 10284 23050
rect 10232 22986 10284 22992
rect 10244 22778 10272 22986
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 9508 22066 9628 22094
rect 9600 22030 9628 22066
rect 9968 22066 10088 22094
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8300 21072 8352 21078
rect 8300 21014 8352 21020
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 8496 20942 8524 21286
rect 8588 21146 8616 21490
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8496 20534 8524 20878
rect 8588 20602 8616 21082
rect 8680 20874 8708 21490
rect 8864 21418 8892 21490
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 8852 21412 8904 21418
rect 8852 21354 8904 21360
rect 8758 21040 8814 21049
rect 8758 20975 8814 20984
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6656 18358 6684 18770
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6656 17814 6684 18294
rect 6748 18086 6776 19110
rect 6932 18970 6960 19110
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18358 7144 18566
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 7116 17678 7144 18294
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 6748 17202 6776 17614
rect 7116 17338 7144 17614
rect 7484 17542 7512 18770
rect 7576 18630 7604 19382
rect 7760 18766 7788 19722
rect 8312 19514 8340 20402
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8022 19272 8078 19281
rect 8022 19207 8078 19216
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7944 18834 7972 19110
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7668 17678 7696 18702
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 18290 7880 18566
rect 8036 18290 8064 19207
rect 8312 18970 8340 19450
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8128 18426 8156 18702
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7852 17202 7880 18022
rect 7944 17882 7972 18158
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 8128 17746 8156 18362
rect 8404 18358 8432 19110
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8496 18290 8524 19926
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6840 16794 6868 17070
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7300 16250 7328 16458
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7392 16114 7420 16934
rect 8220 16590 8248 18158
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1964 13938 1992 14418
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1768 13728 1820 13734
rect 1766 13696 1768 13705
rect 1820 13696 1822 13705
rect 1766 13631 1822 13640
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7002 1624 7346
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1780 6905 1808 7142
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1964 6798 1992 13874
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 8220 13394 8248 16526
rect 8404 15026 8432 17206
rect 8772 16114 8800 20975
rect 9324 20466 9352 21422
rect 9416 21146 9444 21898
rect 9600 21690 9628 21966
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9876 21690 9904 21830
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9692 20874 9720 20946
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9600 19922 9628 20538
rect 9692 20262 9720 20810
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9416 19310 9444 19722
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 8864 18970 8892 19246
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8772 15570 8800 16050
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 8956 12434 8984 15506
rect 9048 15502 9076 17002
rect 9140 16658 9168 17206
rect 9416 16794 9444 19246
rect 9784 17338 9812 20742
rect 9876 20330 9904 21490
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9968 18630 9996 22066
rect 10428 19281 10456 25055
rect 10520 24138 10548 25230
rect 10692 25220 10744 25226
rect 10692 25162 10744 25168
rect 10704 24818 10732 25162
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10980 24886 11008 25094
rect 10968 24880 11020 24886
rect 10968 24822 11020 24828
rect 10692 24812 10744 24818
rect 10612 24772 10692 24800
rect 10612 24614 10640 24772
rect 10692 24754 10744 24760
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10600 24608 10652 24614
rect 10600 24550 10652 24556
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 10704 22642 10732 24618
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11164 22710 11192 23462
rect 11152 22704 11204 22710
rect 11152 22646 11204 22652
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 10612 21146 10640 22442
rect 10704 22030 10732 22578
rect 11152 22500 11204 22506
rect 11152 22442 11204 22448
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22098 11100 22374
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 10692 22024 10744 22030
rect 11164 21978 11192 22442
rect 10692 21966 10744 21972
rect 11072 21962 11192 21978
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11060 21956 11192 21962
rect 11112 21950 11192 21956
rect 11060 21898 11112 21904
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10612 19990 10640 20878
rect 10796 20602 10824 21422
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10414 19272 10470 19281
rect 10414 19207 10470 19216
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9968 17082 9996 18566
rect 10704 18358 10732 20334
rect 10888 19242 10916 21490
rect 11072 21026 11100 21898
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11164 21146 11192 21286
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11072 20998 11192 21026
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10980 20330 11008 20878
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11072 20466 11100 20810
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10980 19360 11008 20266
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11072 20058 11100 20198
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11060 19372 11112 19378
rect 10980 19332 11060 19360
rect 11060 19314 11112 19320
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 11164 19174 11192 20998
rect 11256 20942 11284 21966
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11348 21418 11376 21830
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11256 19310 11284 20878
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11256 18902 11284 19246
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10796 18426 10824 18634
rect 11058 18592 11114 18601
rect 11058 18527 11114 18536
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10704 17814 10732 18294
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 9968 17054 10088 17082
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9968 16590 9996 16934
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9140 14618 9168 14962
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8956 12406 9076 12434
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6564 2650 6592 12310
rect 9048 2922 9076 12406
rect 9232 6914 9260 15438
rect 9324 14550 9352 15846
rect 9956 15496 10008 15502
rect 9954 15464 9956 15473
rect 10008 15464 10010 15473
rect 9954 15399 10010 15408
rect 9968 15162 9996 15399
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10060 14890 10088 17054
rect 10428 16266 10456 17478
rect 10520 17270 10548 17478
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10428 16238 10548 16266
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10336 15978 10364 16050
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10336 15502 10364 15914
rect 10324 15496 10376 15502
rect 10520 15450 10548 16238
rect 10324 15438 10376 15444
rect 10336 15026 10364 15438
rect 10428 15422 10548 15450
rect 10428 15162 10456 15422
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9324 14414 9352 14486
rect 10244 14482 10272 14758
rect 10336 14482 10364 14962
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 10428 14074 10456 15098
rect 10612 15065 10640 17614
rect 11072 17134 11100 18527
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11164 16794 11192 17206
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10796 15638 10824 16186
rect 10980 16182 11008 16390
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10598 15056 10654 15065
rect 10598 14991 10654 15000
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 9876 13938 9904 14010
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 12850 9904 13670
rect 10520 13394 10548 14350
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9968 12986 9996 13194
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10520 12850 10548 13330
rect 10612 12918 10640 14991
rect 10796 14414 10824 15574
rect 10888 15366 10916 16050
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11242 15600 11298 15609
rect 11348 15570 11376 15914
rect 11440 15910 11468 27406
rect 11716 26625 11744 29106
rect 11900 28966 11928 29106
rect 11888 28960 11940 28966
rect 11888 28902 11940 28908
rect 11900 28762 11928 28902
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11808 28014 11836 28358
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 11992 27130 12020 27406
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 12084 27130 12112 27270
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 11702 26616 11758 26625
rect 11702 26551 11758 26560
rect 12176 26466 12204 31350
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 12256 30184 12308 30190
rect 12256 30126 12308 30132
rect 12532 30184 12584 30190
rect 12532 30126 12584 30132
rect 12268 29034 12296 30126
rect 12544 29782 12572 30126
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12532 29776 12584 29782
rect 12452 29724 12532 29730
rect 12452 29718 12584 29724
rect 12452 29702 12572 29718
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12256 29028 12308 29034
rect 12256 28970 12308 28976
rect 12268 28014 12296 28970
rect 12256 28008 12308 28014
rect 12256 27950 12308 27956
rect 12360 27606 12388 29582
rect 12452 29170 12480 29702
rect 12532 29504 12584 29510
rect 12532 29446 12584 29452
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12544 28914 12572 29446
rect 12636 29238 12664 29990
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 12544 28886 12664 28914
rect 12348 27600 12400 27606
rect 12348 27542 12400 27548
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 12268 26586 12296 27338
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12176 26438 12296 26466
rect 12072 26308 12124 26314
rect 12072 26250 12124 26256
rect 12084 25906 12112 26250
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 11900 24818 11928 25162
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11808 22506 11836 24550
rect 11900 23594 11928 24754
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 23866 12204 24074
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 11888 23588 11940 23594
rect 11888 23530 11940 23536
rect 12268 22710 12296 26438
rect 12452 26042 12480 27270
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 11796 22500 11848 22506
rect 11796 22442 11848 22448
rect 11808 21554 11836 22442
rect 12268 22234 12296 22510
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11900 21010 11928 21898
rect 11980 21616 12032 21622
rect 11980 21558 12032 21564
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11532 20602 11560 20946
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11716 20466 11744 20878
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11808 19854 11836 20470
rect 11900 20330 11928 20946
rect 11992 20466 12020 21558
rect 12256 21140 12308 21146
rect 12360 21128 12388 22034
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12452 21146 12480 21966
rect 12544 21690 12572 23666
rect 12636 22030 12664 28886
rect 12728 27538 12756 30738
rect 12808 28484 12860 28490
rect 12808 28426 12860 28432
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 12728 27062 12756 27474
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12728 25226 12756 26998
rect 12716 25220 12768 25226
rect 12716 25162 12768 25168
rect 12728 24818 12756 25162
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12820 23730 12848 28426
rect 12912 28082 12940 32846
rect 13544 32768 13596 32774
rect 13544 32710 13596 32716
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13188 32026 13216 32370
rect 12992 32020 13044 32026
rect 12992 31962 13044 31968
rect 13176 32020 13228 32026
rect 13176 31962 13228 31968
rect 13004 30938 13032 31962
rect 13556 31754 13584 32710
rect 13832 32298 13860 33458
rect 13924 33318 13952 34002
rect 14372 33992 14424 33998
rect 14372 33934 14424 33940
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15936 33992 15988 33998
rect 15936 33934 15988 33940
rect 14004 33856 14056 33862
rect 14004 33798 14056 33804
rect 14016 33454 14044 33798
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 13912 33312 13964 33318
rect 13912 33254 13964 33260
rect 14384 32910 14412 33934
rect 14648 33856 14700 33862
rect 14648 33798 14700 33804
rect 14372 32904 14424 32910
rect 14372 32846 14424 32852
rect 14384 32570 14412 32846
rect 14372 32564 14424 32570
rect 14372 32506 14424 32512
rect 13820 32292 13872 32298
rect 13820 32234 13872 32240
rect 14384 31958 14412 32506
rect 14660 32502 14688 33798
rect 15292 33516 15344 33522
rect 15292 33458 15344 33464
rect 14924 33312 14976 33318
rect 14924 33254 14976 33260
rect 14832 32768 14884 32774
rect 14832 32710 14884 32716
rect 14648 32496 14700 32502
rect 14648 32438 14700 32444
rect 14556 32360 14608 32366
rect 14556 32302 14608 32308
rect 14568 32230 14596 32302
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14372 31952 14424 31958
rect 14372 31894 14424 31900
rect 14188 31884 14240 31890
rect 14188 31826 14240 31832
rect 13464 31726 13584 31754
rect 13728 31748 13780 31754
rect 13268 31408 13320 31414
rect 13268 31350 13320 31356
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 13176 31340 13228 31346
rect 13176 31282 13228 31288
rect 12992 30932 13044 30938
rect 12992 30874 13044 30880
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13004 30190 13032 30670
rect 13096 30598 13124 31282
rect 13188 30841 13216 31282
rect 13174 30832 13230 30841
rect 13174 30767 13230 30776
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 12992 30184 13044 30190
rect 12992 30126 13044 30132
rect 13096 29646 13124 30534
rect 13188 30394 13216 30670
rect 13176 30388 13228 30394
rect 13176 30330 13228 30336
rect 13084 29640 13136 29646
rect 13084 29582 13136 29588
rect 13280 29306 13308 31350
rect 13464 30802 13492 31726
rect 13728 31690 13780 31696
rect 13544 31204 13596 31210
rect 13544 31146 13596 31152
rect 13452 30796 13504 30802
rect 13452 30738 13504 30744
rect 13556 30258 13584 31146
rect 13740 30666 13768 31690
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13544 30252 13596 30258
rect 13544 30194 13596 30200
rect 13636 30184 13688 30190
rect 13636 30126 13688 30132
rect 13544 30116 13596 30122
rect 13544 30058 13596 30064
rect 13268 29300 13320 29306
rect 13268 29242 13320 29248
rect 13556 29238 13584 30058
rect 13648 29714 13676 30126
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13544 29232 13596 29238
rect 13544 29174 13596 29180
rect 12900 28076 12952 28082
rect 12900 28018 12952 28024
rect 13450 27568 13506 27577
rect 13450 27503 13506 27512
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 13096 26586 13124 27406
rect 13268 26784 13320 26790
rect 13268 26726 13320 26732
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 12900 26308 12952 26314
rect 12900 26250 12952 26256
rect 12912 25906 12940 26250
rect 13280 25906 13308 26726
rect 13464 26314 13492 27503
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12820 23322 12848 23666
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22234 12756 22510
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12308 21100 12388 21128
rect 12256 21082 12308 21088
rect 12360 20942 12388 21100
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12544 20942 12572 21422
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12176 20466 12204 20742
rect 11980 20460 12032 20466
rect 12164 20460 12216 20466
rect 12032 20420 12112 20448
rect 11980 20402 12032 20408
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11900 19990 11928 20266
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11992 19854 12020 20266
rect 12084 19854 12112 20420
rect 12164 20402 12216 20408
rect 12820 20346 12848 22442
rect 12820 20318 12940 20346
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12728 19446 12756 19790
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 16250 11560 17682
rect 11716 17542 11744 18022
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11900 17134 11928 18226
rect 12084 17678 12112 18226
rect 12176 18222 12204 18566
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 12176 16658 12204 18158
rect 12452 17202 12480 18838
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12544 17882 12572 18022
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12636 17338 12664 19110
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12728 17338 12756 18226
rect 12820 17882 12848 19314
rect 12912 18766 12940 20318
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 13004 18358 13032 24074
rect 13188 23730 13216 25638
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13372 24750 13400 25434
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13188 20602 13216 23666
rect 13280 23526 13308 24006
rect 13372 23730 13400 24686
rect 13464 24206 13492 25094
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13464 23662 13492 24142
rect 13452 23656 13504 23662
rect 13452 23598 13504 23604
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 19854 13124 20198
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13188 19334 13216 20334
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13280 19514 13308 19790
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13096 19306 13216 19334
rect 13268 19372 13320 19378
rect 13372 19360 13400 19722
rect 13452 19372 13504 19378
rect 13372 19332 13452 19360
rect 13268 19314 13320 19320
rect 13452 19314 13504 19320
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 13004 17542 13032 18022
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 11888 16652 11940 16658
rect 11716 16612 11888 16640
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11716 16114 11744 16612
rect 11888 16594 11940 16600
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11242 15535 11244 15544
rect 11296 15535 11298 15544
rect 11336 15564 11388 15570
rect 11244 15506 11296 15512
rect 11336 15506 11388 15512
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 14618 10916 15302
rect 11716 15026 11744 15846
rect 11808 15570 11836 16458
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12268 16114 12296 16390
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 11900 15706 11928 16050
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 15201 11836 15506
rect 11794 15192 11850 15201
rect 11900 15162 11928 15642
rect 11980 15496 12032 15502
rect 11978 15464 11980 15473
rect 12032 15464 12034 15473
rect 11978 15399 12034 15408
rect 11794 15127 11850 15136
rect 11888 15156 11940 15162
rect 11808 15026 11836 15127
rect 11888 15098 11940 15104
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 12176 14618 12204 15846
rect 12268 15162 12296 16050
rect 12636 15638 12664 16118
rect 12728 16114 12756 16526
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12820 15910 12848 16934
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12820 15434 12848 15846
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10796 12850 10824 13670
rect 10888 12986 10916 13942
rect 11808 13938 11836 14350
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 10980 13530 11008 13874
rect 12360 13870 12388 14758
rect 12544 14618 12572 14962
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12636 13802 12664 14826
rect 12912 14618 12940 16050
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13004 15026 13032 15846
rect 13096 15502 13124 19306
rect 13280 17882 13308 19314
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13096 15026 13124 15438
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12820 14006 12848 14418
rect 13096 14414 13124 14962
rect 13188 14822 13216 17614
rect 13464 16590 13492 19314
rect 13556 18290 13584 29174
rect 13648 27674 13676 29650
rect 13740 29646 13768 30602
rect 14200 30326 14228 31826
rect 14384 31822 14412 31894
rect 14372 31816 14424 31822
rect 14372 31758 14424 31764
rect 14384 31346 14412 31758
rect 14568 31754 14596 32166
rect 14648 31816 14700 31822
rect 14646 31784 14648 31793
rect 14700 31784 14702 31793
rect 14464 31748 14516 31754
rect 14464 31690 14516 31696
rect 14556 31748 14608 31754
rect 14646 31719 14702 31728
rect 14556 31690 14608 31696
rect 14372 31340 14424 31346
rect 14372 31282 14424 31288
rect 14372 31204 14424 31210
rect 14372 31146 14424 31152
rect 14384 30802 14412 31146
rect 14476 31142 14504 31690
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14372 30796 14424 30802
rect 14372 30738 14424 30744
rect 14188 30320 14240 30326
rect 14188 30262 14240 30268
rect 14384 30138 14412 30738
rect 14568 30326 14596 31690
rect 14844 31142 14872 32710
rect 14936 31929 14964 33254
rect 15304 32366 15332 33458
rect 15488 32910 15516 33934
rect 15948 33658 15976 33934
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 15752 33312 15804 33318
rect 15752 33254 15804 33260
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 15384 32836 15436 32842
rect 15384 32778 15436 32784
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 14922 31920 14978 31929
rect 14922 31855 14978 31864
rect 14832 31136 14884 31142
rect 14832 31078 14884 31084
rect 14648 30592 14700 30598
rect 14648 30534 14700 30540
rect 14832 30592 14884 30598
rect 14832 30534 14884 30540
rect 14556 30320 14608 30326
rect 14556 30262 14608 30268
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14476 30138 14504 30194
rect 14384 30110 14504 30138
rect 14384 29850 14412 30110
rect 14464 30048 14516 30054
rect 14464 29990 14516 29996
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 14280 28756 14332 28762
rect 14280 28698 14332 28704
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 13636 27668 13688 27674
rect 13636 27610 13688 27616
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 13648 26994 13676 27474
rect 13728 27464 13780 27470
rect 13728 27406 13780 27412
rect 13740 26994 13768 27406
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 13924 27062 13952 27338
rect 13912 27056 13964 27062
rect 13912 26998 13964 27004
rect 13636 26988 13688 26994
rect 13636 26930 13688 26936
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 13648 25906 13676 26930
rect 13726 26752 13782 26761
rect 13726 26687 13782 26696
rect 13740 26382 13768 26687
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13636 25696 13688 25702
rect 13636 25638 13688 25644
rect 13648 24750 13676 25638
rect 13636 24744 13688 24750
rect 13636 24686 13688 24692
rect 14108 24206 14136 28018
rect 14292 27470 14320 28698
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14292 27130 14320 27270
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14384 26330 14412 29786
rect 14476 29510 14504 29990
rect 14660 29850 14688 30534
rect 14648 29844 14700 29850
rect 14648 29786 14700 29792
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14568 29510 14596 29582
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14556 29504 14608 29510
rect 14556 29446 14608 29452
rect 14476 27062 14504 29446
rect 14660 28694 14688 29786
rect 14740 29776 14792 29782
rect 14740 29718 14792 29724
rect 14752 29646 14780 29718
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14740 29164 14792 29170
rect 14844 29152 14872 30534
rect 14936 29170 14964 31855
rect 15292 31680 15344 31686
rect 15292 31622 15344 31628
rect 15304 30938 15332 31622
rect 15292 30932 15344 30938
rect 15292 30874 15344 30880
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15108 30184 15160 30190
rect 15108 30126 15160 30132
rect 15016 29844 15068 29850
rect 15016 29786 15068 29792
rect 14792 29124 14872 29152
rect 14924 29164 14976 29170
rect 14740 29106 14792 29112
rect 14924 29106 14976 29112
rect 15028 28994 15056 29786
rect 14936 28966 15056 28994
rect 14648 28688 14700 28694
rect 14648 28630 14700 28636
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14568 27606 14596 28494
rect 14648 28416 14700 28422
rect 14648 28358 14700 28364
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14464 27056 14516 27062
rect 14464 26998 14516 27004
rect 14476 26450 14504 26998
rect 14568 26586 14596 27270
rect 14660 26761 14688 28358
rect 14752 28150 14780 28562
rect 14740 28144 14792 28150
rect 14740 28086 14792 28092
rect 14832 27464 14884 27470
rect 14830 27432 14832 27441
rect 14936 27452 14964 28966
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 15028 27606 15056 28494
rect 15016 27600 15068 27606
rect 15016 27542 15068 27548
rect 14884 27432 14964 27452
rect 14886 27424 14964 27432
rect 15016 27464 15068 27470
rect 15016 27406 15068 27412
rect 14830 27367 14886 27376
rect 14844 26790 14872 27367
rect 14922 27024 14978 27033
rect 14922 26959 14978 26968
rect 14832 26784 14884 26790
rect 14646 26752 14702 26761
rect 14832 26726 14884 26732
rect 14646 26687 14702 26696
rect 14936 26586 14964 26959
rect 14556 26580 14608 26586
rect 14556 26522 14608 26528
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 14464 26444 14516 26450
rect 14516 26404 14688 26432
rect 14464 26386 14516 26392
rect 14384 26302 14504 26330
rect 14372 25696 14424 25702
rect 14372 25638 14424 25644
rect 14384 25226 14412 25638
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14384 24886 14412 25162
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14108 23594 14136 24142
rect 14200 23866 14228 24346
rect 14278 23896 14334 23905
rect 14188 23860 14240 23866
rect 14278 23831 14280 23840
rect 14188 23802 14240 23808
rect 14332 23831 14334 23840
rect 14280 23802 14332 23808
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 14096 23588 14148 23594
rect 14096 23530 14148 23536
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13648 21690 13676 21966
rect 13924 21962 13952 23530
rect 14476 22982 14504 26302
rect 14556 26308 14608 26314
rect 14556 26250 14608 26256
rect 14568 25294 14596 26250
rect 14660 25702 14688 26404
rect 14738 26344 14794 26353
rect 14738 26279 14794 26288
rect 14648 25696 14700 25702
rect 14648 25638 14700 25644
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14568 24818 14596 25230
rect 14752 24818 14780 26279
rect 15028 25906 15056 27406
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14292 22030 14320 22442
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 13912 21956 13964 21962
rect 13912 21898 13964 21904
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 14278 20496 14334 20505
rect 14278 20431 14280 20440
rect 14332 20431 14334 20440
rect 14280 20402 14332 20408
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14476 20233 14504 20334
rect 14568 20262 14596 24754
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14660 20398 14688 20946
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14556 20256 14608 20262
rect 14462 20224 14518 20233
rect 14556 20198 14608 20204
rect 14462 20159 14518 20168
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13740 19310 13768 19790
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13832 19378 13860 19722
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13648 18970 13676 19110
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13556 17678 13584 18226
rect 13648 17814 13676 18634
rect 13740 17882 13768 19246
rect 13912 19168 13964 19174
rect 13832 19128 13912 19156
rect 13832 18290 13860 19128
rect 13912 19110 13964 19116
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18426 13952 18566
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14016 18290 14044 18634
rect 14108 18426 14136 18702
rect 14292 18698 14320 19654
rect 14476 19378 14504 20159
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14568 18766 14596 20198
rect 14752 19922 14780 20538
rect 14844 20466 14872 25842
rect 14924 25152 14976 25158
rect 14922 25120 14924 25129
rect 14976 25120 14978 25129
rect 14922 25055 14978 25064
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 14936 23866 14964 24074
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14922 23760 14978 23769
rect 14922 23695 14978 23704
rect 14936 20584 14964 23695
rect 15120 23118 15148 30126
rect 15304 30054 15332 30602
rect 15292 30048 15344 30054
rect 15292 29990 15344 29996
rect 15304 29782 15332 29990
rect 15292 29776 15344 29782
rect 15292 29718 15344 29724
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15304 29306 15332 29582
rect 15292 29300 15344 29306
rect 15292 29242 15344 29248
rect 15396 28558 15424 32778
rect 15488 32774 15516 32846
rect 15476 32768 15528 32774
rect 15476 32710 15528 32716
rect 15488 32434 15516 32710
rect 15580 32502 15608 32914
rect 15568 32496 15620 32502
rect 15764 32450 15792 33254
rect 16132 32910 16160 33798
rect 16224 33454 16252 34002
rect 16212 33448 16264 33454
rect 16210 33416 16212 33425
rect 16264 33416 16266 33425
rect 16210 33351 16266 33360
rect 17040 33380 17092 33386
rect 17040 33322 17092 33328
rect 16488 33312 16540 33318
rect 16488 33254 16540 33260
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 16040 32570 16068 32710
rect 16028 32564 16080 32570
rect 16028 32506 16080 32512
rect 15568 32438 15620 32444
rect 15476 32428 15528 32434
rect 15476 32370 15528 32376
rect 15488 31890 15516 32370
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15580 31872 15608 32438
rect 15672 32434 15792 32450
rect 16500 32434 16528 33254
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 15660 32428 15792 32434
rect 15712 32422 15792 32428
rect 15660 32370 15712 32376
rect 15660 31884 15712 31890
rect 15580 31844 15660 31872
rect 15476 31748 15528 31754
rect 15476 31690 15528 31696
rect 15488 29850 15516 31690
rect 15580 30190 15608 31844
rect 15660 31826 15712 31832
rect 15764 30938 15792 32422
rect 15844 32428 15896 32434
rect 16488 32428 16540 32434
rect 15896 32388 15976 32416
rect 15844 32370 15896 32376
rect 15948 31958 15976 32388
rect 16488 32370 16540 32376
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 15936 31952 15988 31958
rect 15842 31920 15898 31929
rect 15936 31894 15988 31900
rect 15842 31855 15844 31864
rect 15896 31855 15898 31864
rect 15844 31826 15896 31832
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 15752 30932 15804 30938
rect 15752 30874 15804 30880
rect 15651 30660 15703 30666
rect 15651 30602 15703 30608
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15672 29578 15700 30602
rect 15764 30258 15792 30874
rect 15844 30864 15896 30870
rect 15844 30806 15896 30812
rect 15752 30252 15804 30258
rect 15752 30194 15804 30200
rect 15856 30122 15884 30806
rect 16040 30734 16068 31078
rect 16224 30938 16252 32166
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16212 30932 16264 30938
rect 16212 30874 16264 30880
rect 16028 30728 16080 30734
rect 16028 30670 16080 30676
rect 16316 30394 16344 31282
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 15764 29646 15792 29990
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15660 29572 15712 29578
rect 15660 29514 15712 29520
rect 15764 29238 15792 29582
rect 15752 29232 15804 29238
rect 15752 29174 15804 29180
rect 15764 28994 15792 29174
rect 15672 28966 15792 28994
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15212 27606 15240 28426
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15200 27600 15252 27606
rect 15200 27542 15252 27548
rect 15200 26988 15252 26994
rect 15304 26976 15332 28358
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15476 27940 15528 27946
rect 15476 27882 15528 27888
rect 15488 27470 15516 27882
rect 15580 27538 15608 27950
rect 15568 27532 15620 27538
rect 15568 27474 15620 27480
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15384 27328 15436 27334
rect 15384 27270 15436 27276
rect 15252 26948 15332 26976
rect 15200 26930 15252 26936
rect 15212 26042 15240 26930
rect 15396 26382 15424 27270
rect 15488 26994 15516 27406
rect 15568 27124 15620 27130
rect 15568 27066 15620 27072
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15476 26784 15528 26790
rect 15474 26752 15476 26761
rect 15528 26752 15530 26761
rect 15474 26687 15530 26696
rect 15580 26586 15608 27066
rect 15672 26926 15700 28966
rect 15660 26920 15712 26926
rect 15660 26862 15712 26868
rect 15856 26586 15884 30058
rect 16040 29850 16068 30262
rect 16684 30258 16712 33050
rect 16764 32768 16816 32774
rect 16764 32710 16816 32716
rect 16776 32298 16804 32710
rect 16764 32292 16816 32298
rect 16764 32234 16816 32240
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16488 30048 16540 30054
rect 16488 29990 16540 29996
rect 16500 29850 16528 29990
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16500 29753 16528 29786
rect 16486 29744 16542 29753
rect 16486 29679 16542 29688
rect 16488 29640 16540 29646
rect 16488 29582 16540 29588
rect 16304 29504 16356 29510
rect 16304 29446 16356 29452
rect 16212 29300 16264 29306
rect 16212 29242 16264 29248
rect 16224 27878 16252 29242
rect 16212 27872 16264 27878
rect 16212 27814 16264 27820
rect 16224 27690 16252 27814
rect 16132 27662 16252 27690
rect 16132 27470 16160 27662
rect 16212 27600 16264 27606
rect 16210 27568 16212 27577
rect 16264 27568 16266 27577
rect 16210 27503 16266 27512
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 16132 26926 16160 27406
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 16316 26738 16344 29446
rect 16396 28416 16448 28422
rect 16396 28358 16448 28364
rect 16408 28014 16436 28358
rect 16396 28008 16448 28014
rect 16396 27950 16448 27956
rect 16408 26858 16436 27950
rect 16500 26994 16528 29582
rect 16776 29170 16804 32234
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16960 30258 16988 31078
rect 17052 30734 17080 33322
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17236 30938 17264 32370
rect 17328 31346 17356 34070
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 18052 32836 18104 32842
rect 18052 32778 18104 32784
rect 17684 32224 17736 32230
rect 17684 32166 17736 32172
rect 17696 31822 17724 32166
rect 18064 31958 18092 32778
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 27172 32026 27200 37198
rect 32876 37126 32904 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 32956 37256 33008 37262
rect 32956 37198 33008 37204
rect 37832 37256 37884 37262
rect 37832 37198 37884 37204
rect 32864 37120 32916 37126
rect 32864 37062 32916 37068
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 18052 31952 18104 31958
rect 18052 31894 18104 31900
rect 17684 31816 17736 31822
rect 17684 31758 17736 31764
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 17316 31340 17368 31346
rect 17316 31282 17368 31288
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16764 29164 16816 29170
rect 16764 29106 16816 29112
rect 16776 28626 16804 29106
rect 17052 28762 17080 30670
rect 17328 30326 17356 31282
rect 17880 30938 17908 31282
rect 18972 31272 19024 31278
rect 18892 31220 18972 31226
rect 18892 31214 19024 31220
rect 18892 31198 19012 31214
rect 18892 31142 18920 31198
rect 18880 31136 18932 31142
rect 18880 31078 18932 31084
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 17316 30320 17368 30326
rect 17316 30262 17368 30268
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17144 29170 17172 29990
rect 18432 29850 18460 30670
rect 18696 30592 18748 30598
rect 18696 30534 18748 30540
rect 18708 30394 18736 30534
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 17880 29306 17908 29446
rect 17868 29300 17920 29306
rect 17868 29242 17920 29248
rect 17592 29232 17644 29238
rect 17592 29174 17644 29180
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 17040 28756 17092 28762
rect 17040 28698 17092 28704
rect 17144 28642 17172 29106
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16764 28620 16816 28626
rect 16764 28562 16816 28568
rect 17052 28614 17172 28642
rect 16592 27674 16620 28562
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 16488 26988 16540 26994
rect 16488 26930 16540 26936
rect 16868 26858 16896 28018
rect 16948 27872 17000 27878
rect 16948 27814 17000 27820
rect 16960 27402 16988 27814
rect 17052 27538 17080 28614
rect 17224 28416 17276 28422
rect 17224 28358 17276 28364
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16948 27396 17000 27402
rect 16948 27338 17000 27344
rect 16948 26988 17000 26994
rect 17052 26976 17080 27474
rect 17144 27334 17172 28018
rect 17236 27538 17264 28358
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17000 26948 17080 26976
rect 16948 26930 17000 26936
rect 16396 26852 16448 26858
rect 16396 26794 16448 26800
rect 16856 26852 16908 26858
rect 16856 26794 16908 26800
rect 16960 26738 16988 26930
rect 17144 26761 17172 27270
rect 17420 27130 17448 27814
rect 17604 27402 17632 29174
rect 18236 29164 18288 29170
rect 18236 29106 18288 29112
rect 17960 29096 18012 29102
rect 17958 29064 17960 29073
rect 18012 29064 18014 29073
rect 17958 28999 18014 29008
rect 18248 28966 18276 29106
rect 18236 28960 18288 28966
rect 18236 28902 18288 28908
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 18788 28688 18840 28694
rect 18788 28630 18840 28636
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17972 27470 18000 28494
rect 18144 28484 18196 28490
rect 18144 28426 18196 28432
rect 18156 28082 18184 28426
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 18156 27470 18184 28018
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17972 27130 18000 27406
rect 17408 27124 17460 27130
rect 17408 27066 17460 27072
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 15568 26580 15620 26586
rect 15568 26522 15620 26528
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15384 26376 15436 26382
rect 15384 26318 15436 26324
rect 15200 26036 15252 26042
rect 15200 25978 15252 25984
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15304 24800 15332 25638
rect 15396 25158 15424 26318
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15764 24954 15792 25842
rect 15856 25498 15884 26522
rect 15948 26382 15976 26726
rect 16132 26450 16160 26726
rect 16316 26710 16436 26738
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 16026 26344 16082 26353
rect 16026 26279 16028 26288
rect 16080 26279 16082 26288
rect 16028 26250 16080 26256
rect 16040 25974 16068 26250
rect 16028 25968 16080 25974
rect 16028 25910 16080 25916
rect 15844 25492 15896 25498
rect 15844 25434 15896 25440
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15384 24812 15436 24818
rect 15304 24772 15384 24800
rect 15384 24754 15436 24760
rect 15396 24721 15424 24754
rect 15382 24712 15438 24721
rect 15382 24647 15438 24656
rect 15658 24168 15714 24177
rect 15658 24103 15714 24112
rect 15672 24070 15700 24103
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 15120 20806 15148 22918
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15212 21554 15240 21830
rect 15304 21706 15332 22510
rect 15396 22030 15424 23122
rect 15856 22982 15884 25434
rect 16040 25294 16068 25910
rect 16120 25356 16172 25362
rect 16120 25298 16172 25304
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 16132 24818 16160 25298
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24993 16252 25094
rect 16210 24984 16266 24993
rect 16210 24919 16266 24928
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 16040 23322 16068 23666
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 16132 23202 16160 24754
rect 16408 24206 16436 26710
rect 16868 26710 16988 26738
rect 17130 26752 17186 26761
rect 16670 26616 16726 26625
rect 16670 26551 16726 26560
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16212 23860 16264 23866
rect 16212 23802 16264 23808
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 16040 23174 16160 23202
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15304 21678 15516 21706
rect 15488 21622 15516 21678
rect 15476 21616 15528 21622
rect 15476 21558 15528 21564
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 14936 20556 15148 20584
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14844 19514 14872 20402
rect 15014 20360 15070 20369
rect 14924 20324 14976 20330
rect 15014 20295 15070 20304
rect 14924 20266 14976 20272
rect 14936 19990 14964 20266
rect 14924 19984 14976 19990
rect 14924 19926 14976 19932
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13648 16998 13676 17750
rect 13832 17678 13860 18226
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14108 17746 14136 18158
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 14476 17202 14504 17750
rect 15028 17678 15056 20295
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15028 17202 15056 17274
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15120 17066 15148 20556
rect 15212 19854 15240 21490
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15304 21146 15332 21286
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15304 18834 15332 19246
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 15212 16726 15240 18226
rect 15396 18222 15424 21286
rect 15488 18970 15516 21558
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15580 18358 15608 22714
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15672 21690 15700 22646
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 15752 22432 15804 22438
rect 15752 22374 15804 22380
rect 15764 21962 15792 22374
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15672 20942 15700 21626
rect 15856 21146 15884 22510
rect 15948 21962 15976 23122
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15856 20942 15884 21082
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15948 20874 15976 21898
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15672 20262 15700 20402
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15764 20058 15792 20402
rect 15856 20346 15884 20470
rect 15948 20466 15976 20538
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15856 20318 15976 20346
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15658 19544 15714 19553
rect 15764 19514 15792 19994
rect 15658 19479 15660 19488
rect 15712 19479 15714 19488
rect 15752 19508 15804 19514
rect 15660 19450 15712 19456
rect 15752 19450 15804 19456
rect 15856 19446 15884 20198
rect 15948 19922 15976 20318
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 16040 19854 16068 23174
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16132 19514 16160 22918
rect 16224 19718 16252 23802
rect 16316 23730 16344 24006
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16316 23633 16344 23666
rect 16302 23624 16358 23633
rect 16302 23559 16358 23568
rect 16408 23118 16436 24142
rect 16500 23866 16528 25298
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 16592 23186 16620 24142
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16592 22778 16620 22986
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16316 20330 16344 20402
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16316 19836 16344 19926
rect 16316 19808 16436 19836
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16316 19553 16344 19654
rect 16302 19544 16358 19553
rect 16120 19508 16172 19514
rect 16302 19479 16358 19488
rect 16120 19450 16172 19456
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15304 17882 15332 18158
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15304 17202 15332 17614
rect 15488 17610 15516 17818
rect 16316 17678 16344 18838
rect 16408 18834 16436 19808
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16500 18714 16528 21966
rect 16592 18902 16620 22714
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16408 18686 16528 18714
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17202 15700 17478
rect 16132 17338 16160 17614
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15304 16946 15332 17138
rect 15304 16918 15424 16946
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13556 16046 13584 16458
rect 15304 16114 15332 16730
rect 15396 16250 15424 16918
rect 15566 16688 15622 16697
rect 15566 16623 15568 16632
rect 15620 16623 15622 16632
rect 15568 16594 15620 16600
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15488 16182 15516 16458
rect 15672 16454 15700 17138
rect 15764 16590 15792 17138
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13556 15570 13584 15982
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14482 13216 14758
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11624 13326 11652 13670
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 12820 12782 12848 13942
rect 13188 13938 13216 14214
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13280 12850 13308 15302
rect 13556 15026 13584 15506
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13464 12986 13492 14350
rect 13556 13938 13584 14418
rect 13740 14414 13768 14894
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13530 13584 13874
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13556 12850 13584 13466
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 13740 12714 13768 14350
rect 13832 13938 13860 14758
rect 13924 14618 13952 15846
rect 14278 15192 14334 15201
rect 14278 15127 14334 15136
rect 14292 15026 14320 15127
rect 14568 15065 14596 15846
rect 15120 15162 15148 16050
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15638 15424 15982
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15384 15496 15436 15502
rect 15488 15450 15516 16118
rect 15436 15444 15516 15450
rect 15384 15438 15516 15444
rect 15396 15422 15516 15438
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 14554 15056 14610 15065
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14464 15020 14516 15026
rect 14554 14991 14556 15000
rect 14464 14962 14516 14968
rect 14608 14991 14610 15000
rect 14556 14962 14608 14968
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14016 14550 14044 14758
rect 14476 14618 14504 14962
rect 15212 14958 15240 15302
rect 15396 14958 15424 15422
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 14384 13530 14412 14350
rect 15028 14074 15056 14350
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 15028 13326 15056 14010
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14752 12986 14780 13194
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 15028 12850 15056 13262
rect 15212 13258 15240 14894
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15304 14414 15332 14826
rect 15396 14822 15424 14894
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15580 14618 15608 16186
rect 15672 15502 15700 16390
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15764 15162 15792 16526
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15856 14958 15884 16050
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15580 14090 15608 14554
rect 15488 14074 15608 14090
rect 15488 14068 15620 14074
rect 15488 14062 15568 14068
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15304 12918 15332 13874
rect 15488 12986 15516 14062
rect 15568 14010 15620 14016
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 9140 6886 9260 6914
rect 9140 3126 9168 6886
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 15304 2514 15332 12854
rect 15580 12850 15608 13874
rect 15948 13326 15976 16934
rect 16040 15910 16068 16934
rect 16132 16794 16160 17274
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16408 16674 16436 18686
rect 16488 18624 16540 18630
rect 16684 18578 16712 26551
rect 16868 25702 16896 26710
rect 17130 26687 17186 26696
rect 17038 26616 17094 26625
rect 17038 26551 17094 26560
rect 17052 26518 17080 26551
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 17144 26296 17172 26687
rect 17052 26268 17172 26296
rect 17316 26308 17368 26314
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16776 23905 16804 24006
rect 16762 23896 16818 23905
rect 16762 23831 16818 23840
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16776 22778 16804 23054
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 21010 16804 21286
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16776 19922 16804 20946
rect 16868 20505 16896 25638
rect 17052 22030 17080 26268
rect 17316 26250 17368 26256
rect 17328 25906 17356 26250
rect 17316 25900 17368 25906
rect 17316 25842 17368 25848
rect 17328 25294 17356 25842
rect 17420 25362 17448 27066
rect 17684 26852 17736 26858
rect 17684 26794 17736 26800
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17408 25356 17460 25362
rect 17408 25298 17460 25304
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 17144 22778 17172 22986
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16854 20496 16910 20505
rect 16854 20431 16910 20440
rect 16960 19922 16988 21490
rect 17052 21486 17080 21830
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16960 18970 16988 19858
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16540 18572 16712 18578
rect 16488 18566 16712 18572
rect 16500 18550 16712 18566
rect 16684 17202 16712 18550
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16868 17134 16896 17682
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16316 16646 16436 16674
rect 16316 16250 16344 16646
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16224 15706 16252 15982
rect 16408 15910 16436 16526
rect 16500 16182 16528 16526
rect 16488 16176 16540 16182
rect 16868 16164 16896 17070
rect 16960 16266 16988 18906
rect 17132 18624 17184 18630
rect 17130 18592 17132 18601
rect 17184 18592 17186 18601
rect 17130 18527 17186 18536
rect 17236 16590 17264 22034
rect 17328 19174 17356 25094
rect 17512 24818 17540 26726
rect 17696 25702 17724 26794
rect 17972 26568 18000 27066
rect 18156 26926 18184 27406
rect 18248 27334 18276 27406
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 18052 26580 18104 26586
rect 17972 26540 18052 26568
rect 18052 26522 18104 26528
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17696 24818 17724 25638
rect 17868 25424 17920 25430
rect 17868 25366 17920 25372
rect 17880 24818 17908 25366
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17972 24886 18000 25094
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17420 22778 17448 23122
rect 17512 23118 17540 24142
rect 17590 23624 17646 23633
rect 17590 23559 17646 23568
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17420 22642 17448 22714
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17512 22166 17540 23054
rect 17604 22642 17632 23559
rect 17972 22982 18000 24822
rect 18064 23338 18092 26522
rect 18156 25974 18184 26862
rect 18248 26382 18276 26930
rect 18340 26586 18368 28630
rect 18696 28212 18748 28218
rect 18696 28154 18748 28160
rect 18512 27940 18564 27946
rect 18512 27882 18564 27888
rect 18524 27674 18552 27882
rect 18708 27674 18736 28154
rect 18800 27878 18828 28630
rect 18788 27872 18840 27878
rect 18788 27814 18840 27820
rect 18512 27668 18564 27674
rect 18512 27610 18564 27616
rect 18696 27668 18748 27674
rect 18696 27610 18748 27616
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18432 27062 18460 27270
rect 18420 27056 18472 27062
rect 18420 26998 18472 27004
rect 18420 26852 18472 26858
rect 18420 26794 18472 26800
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18432 26382 18460 26794
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 18248 23866 18276 26318
rect 18524 25362 18552 27610
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 18616 25974 18644 27542
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18616 25242 18644 25910
rect 18708 25412 18736 27610
rect 18892 26926 18920 31078
rect 19248 30660 19300 30666
rect 19248 30602 19300 30608
rect 19340 30660 19392 30666
rect 19340 30602 19392 30608
rect 19064 30592 19116 30598
rect 19064 30534 19116 30540
rect 19076 30258 19104 30534
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 19076 29220 19104 30194
rect 19156 29232 19208 29238
rect 19076 29192 19156 29220
rect 19076 28694 19104 29192
rect 19156 29174 19208 29180
rect 19064 28688 19116 28694
rect 19064 28630 19116 28636
rect 18972 28552 19024 28558
rect 19260 28540 19288 30602
rect 19352 30190 19380 30602
rect 19340 30184 19392 30190
rect 19340 30126 19392 30132
rect 19352 29714 19380 30126
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19352 29034 19380 29650
rect 19444 29102 19472 31078
rect 19996 30870 20024 31758
rect 20076 31680 20128 31686
rect 20076 31622 20128 31628
rect 20088 31414 20116 31622
rect 20076 31408 20128 31414
rect 20076 31350 20128 31356
rect 25320 31408 25372 31414
rect 25320 31350 25372 31356
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 23112 31340 23164 31346
rect 23112 31282 23164 31288
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 22020 31142 22048 31282
rect 23020 31204 23072 31210
rect 23020 31146 23072 31152
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 22284 31136 22336 31142
rect 22284 31078 22336 31084
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 20916 30802 20944 31078
rect 20904 30796 20956 30802
rect 20904 30738 20956 30744
rect 21180 30796 21232 30802
rect 21180 30738 21232 30744
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20352 30592 20404 30598
rect 20352 30534 20404 30540
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 20364 30258 20392 30534
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20456 29850 20484 30670
rect 21192 29850 21220 30738
rect 22020 30326 22048 31078
rect 22008 30320 22060 30326
rect 22008 30262 22060 30268
rect 22296 30122 22324 31078
rect 23032 30802 23060 31146
rect 23020 30796 23072 30802
rect 23020 30738 23072 30744
rect 22560 30728 22612 30734
rect 22560 30670 22612 30676
rect 22572 30258 22600 30670
rect 22560 30252 22612 30258
rect 22560 30194 22612 30200
rect 22284 30116 22336 30122
rect 22284 30058 22336 30064
rect 21456 30048 21508 30054
rect 21456 29990 21508 29996
rect 20444 29844 20496 29850
rect 20444 29786 20496 29792
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 21468 29578 21496 29990
rect 21456 29572 21508 29578
rect 21456 29514 21508 29520
rect 20076 29504 20128 29510
rect 20076 29446 20128 29452
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 20088 29306 20116 29446
rect 20076 29300 20128 29306
rect 20076 29242 20128 29248
rect 20548 29170 20576 29446
rect 21468 29170 21496 29514
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19340 29028 19392 29034
rect 19340 28970 19392 28976
rect 18972 28494 19024 28500
rect 19076 28512 19288 28540
rect 18984 28218 19012 28494
rect 18972 28212 19024 28218
rect 18972 28154 19024 28160
rect 18972 26988 19024 26994
rect 18972 26930 19024 26936
rect 18880 26920 18932 26926
rect 18880 26862 18932 26868
rect 18892 26586 18920 26862
rect 18880 26580 18932 26586
rect 18880 26522 18932 26528
rect 18984 26042 19012 26930
rect 18972 26036 19024 26042
rect 18972 25978 19024 25984
rect 18880 25424 18932 25430
rect 18708 25384 18828 25412
rect 18616 25214 18736 25242
rect 18708 25158 18736 25214
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18800 24800 18828 25384
rect 18880 25366 18932 25372
rect 18892 25294 18920 25366
rect 18880 25288 18932 25294
rect 18932 25248 19012 25276
rect 18880 25230 18932 25236
rect 18880 25152 18932 25158
rect 18880 25094 18932 25100
rect 18892 24954 18920 25094
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18432 24772 18828 24800
rect 18880 24812 18932 24818
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18064 23322 18184 23338
rect 18064 23316 18196 23322
rect 18064 23310 18144 23316
rect 18144 23258 18196 23264
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 17500 22160 17552 22166
rect 17500 22102 17552 22108
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17420 21690 17448 21830
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17512 20806 17540 21014
rect 17604 20874 17632 21966
rect 17880 21690 17908 22034
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17696 21146 17724 21490
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17880 20942 17908 21626
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17592 20868 17644 20874
rect 17592 20810 17644 20816
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17788 20233 17816 20402
rect 17880 20262 17908 20878
rect 18052 20324 18104 20330
rect 18052 20266 18104 20272
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 17868 20256 17920 20262
rect 17774 20224 17830 20233
rect 17868 20198 17920 20204
rect 17774 20159 17830 20168
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17604 18698 17632 19246
rect 17696 18970 17724 19722
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17788 18970 17816 19314
rect 17880 19310 17908 19722
rect 18064 19514 18092 20266
rect 18156 20058 18184 20266
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18156 19514 18184 19994
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17788 18766 17816 18906
rect 17972 18766 18000 19110
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 18064 18714 18092 19450
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18156 18902 18184 19314
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18144 18760 18196 18766
rect 18064 18708 18144 18714
rect 18064 18702 18196 18708
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17592 18692 17644 18698
rect 18064 18686 18184 18702
rect 17592 18634 17644 18640
rect 17512 18290 17540 18634
rect 17776 18352 17828 18358
rect 17776 18294 17828 18300
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 17202 17540 18226
rect 17788 17882 17816 18294
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17972 17882 18000 18090
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 16960 16238 17172 16266
rect 17040 16176 17092 16182
rect 16868 16136 17040 16164
rect 16488 16118 16540 16124
rect 17040 16118 17092 16124
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16316 15570 16344 15846
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16408 15026 16436 15846
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16592 15094 16620 15574
rect 16960 15502 16988 15846
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16500 14278 16528 14962
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 16500 12782 16528 14214
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16592 12714 16620 15030
rect 16776 14890 16804 15438
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 13938 16988 14350
rect 17052 14006 17080 16118
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 17144 13938 17172 16238
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17236 15706 17264 16050
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17236 13938 17264 15370
rect 17328 14550 17356 16390
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17420 15502 17448 16118
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17316 14544 17368 14550
rect 17316 14486 17368 14492
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 16960 13530 16988 13874
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17144 13258 17172 13874
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 17052 12306 17080 12650
rect 17512 12442 17540 17138
rect 18156 17066 18184 17818
rect 18248 17814 18276 22578
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18340 20806 18368 20878
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18326 20224 18382 20233
rect 18326 20159 18382 20168
rect 18340 20058 18368 20159
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18432 19718 18460 24772
rect 18880 24754 18932 24760
rect 18788 24676 18840 24682
rect 18892 24664 18920 24754
rect 18840 24636 18920 24664
rect 18788 24618 18840 24624
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18616 22642 18644 23258
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18708 22506 18736 23598
rect 18984 22778 19012 25248
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18524 21078 18552 21966
rect 18708 21146 18736 21966
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18512 21072 18564 21078
rect 18512 21014 18564 21020
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18340 17354 18368 18362
rect 18420 17604 18472 17610
rect 18420 17546 18472 17552
rect 18248 17326 18368 17354
rect 18432 17338 18460 17546
rect 18420 17332 18472 17338
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17604 16250 17632 16458
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17696 15026 17724 15642
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17696 14618 17724 14962
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17788 14822 17816 14894
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17788 14414 17816 14758
rect 17972 14618 18000 15370
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18064 14482 18092 16594
rect 18248 14890 18276 17326
rect 18420 17274 18472 17280
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18340 16794 18368 17138
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18432 16182 18460 17070
rect 18524 16726 18552 21014
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 19922 18644 20198
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18708 19378 18736 20538
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18984 19310 19012 20946
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18984 19174 19012 19246
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18616 18290 18644 18702
rect 19076 18358 19104 28512
rect 19444 28490 19472 29038
rect 20548 29034 20576 29106
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20916 28694 20944 29106
rect 20996 28960 21048 28966
rect 20996 28902 21048 28908
rect 20904 28688 20956 28694
rect 20904 28630 20956 28636
rect 20720 28620 20772 28626
rect 20720 28562 20772 28568
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 20536 28076 20588 28082
rect 20536 28018 20588 28024
rect 19352 27402 19380 28018
rect 20548 27606 20576 28018
rect 20732 27606 20760 28562
rect 21008 28150 21036 28902
rect 20996 28144 21048 28150
rect 20996 28086 21048 28092
rect 21192 27878 21220 29106
rect 21468 28082 21496 29106
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21180 27872 21232 27878
rect 21180 27814 21232 27820
rect 21272 27872 21324 27878
rect 21272 27814 21324 27820
rect 21284 27674 21312 27814
rect 21272 27668 21324 27674
rect 21272 27610 21324 27616
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 20536 27600 20588 27606
rect 20536 27542 20588 27548
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 19352 27130 19380 27338
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19352 26450 19380 27066
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19260 25974 19288 26182
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 19444 25922 19472 27542
rect 21560 27538 21588 29446
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22112 28082 22140 29106
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22204 28218 22232 28494
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 21548 27532 21600 27538
rect 21548 27474 21600 27480
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19892 26852 19944 26858
rect 19892 26794 19944 26800
rect 19904 26382 19932 26794
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 19892 26376 19944 26382
rect 19944 26336 20024 26364
rect 19892 26318 19944 26324
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19168 25498 19196 25842
rect 19156 25492 19208 25498
rect 19156 25434 19208 25440
rect 19260 24818 19288 25910
rect 19444 25894 19564 25922
rect 19536 25838 19564 25894
rect 19892 25900 19944 25906
rect 19892 25842 19944 25848
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19708 25832 19760 25838
rect 19708 25774 19760 25780
rect 19340 25424 19392 25430
rect 19338 25392 19340 25401
rect 19392 25392 19394 25401
rect 19720 25344 19748 25774
rect 19338 25327 19394 25336
rect 19628 25316 19748 25344
rect 19340 25220 19392 25226
rect 19628 25208 19656 25316
rect 19392 25180 19656 25208
rect 19706 25256 19762 25265
rect 19706 25191 19708 25200
rect 19340 25162 19392 25168
rect 19760 25191 19762 25200
rect 19708 25162 19760 25168
rect 19904 25140 19932 25842
rect 19996 25838 20024 26336
rect 20088 25906 20116 26386
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19996 25294 20024 25774
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19338 25120 19394 25129
rect 19904 25112 20024 25140
rect 19338 25055 19394 25064
rect 19352 24954 19380 25055
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19154 24712 19210 24721
rect 19154 24647 19210 24656
rect 19168 24614 19196 24647
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 19168 23662 19196 24210
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19168 18986 19196 23598
rect 19260 22710 19288 24754
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19800 24744 19852 24750
rect 19996 24732 20024 25112
rect 20088 24886 20116 25638
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19852 24704 20024 24732
rect 19800 24686 19852 24692
rect 19352 24290 19380 24686
rect 19708 24676 19760 24682
rect 19708 24618 19760 24624
rect 19720 24410 19748 24618
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19352 24262 19472 24290
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19352 23662 19380 24074
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19352 23186 19380 23598
rect 19444 23322 19472 24262
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19444 22642 19472 22986
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19444 21622 19472 22578
rect 19996 22574 20024 24704
rect 20180 24682 20208 25910
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 20272 24954 20300 25842
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 20088 22982 20116 24278
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 20180 22094 20208 24618
rect 20364 24206 20392 26386
rect 20456 26042 20484 27474
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 22100 27328 22152 27334
rect 22100 27270 22152 27276
rect 20536 26512 20588 26518
rect 20536 26454 20588 26460
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20456 24410 20484 25978
rect 20548 25498 20576 26454
rect 21008 26382 21036 27270
rect 22112 26994 22140 27270
rect 22296 27146 22324 30058
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22388 28558 22416 28902
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22296 27118 22416 27146
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22284 26852 22336 26858
rect 22284 26794 22336 26800
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22100 26512 22152 26518
rect 22100 26454 22152 26460
rect 20996 26376 21048 26382
rect 20996 26318 21048 26324
rect 21732 26240 21784 26246
rect 21732 26182 21784 26188
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20536 25492 20588 25498
rect 20536 25434 20588 25440
rect 20536 24812 20588 24818
rect 20640 24800 20668 25774
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20732 24954 20760 25094
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 20588 24772 20668 24800
rect 20536 24754 20588 24760
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20272 22642 20300 22986
rect 20364 22710 20392 24142
rect 20456 23186 20484 24346
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 20548 23730 20576 24142
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20180 22066 20300 22094
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19628 21078 19656 21490
rect 19996 21486 20024 21966
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20180 21622 20208 21830
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19616 21072 19668 21078
rect 19616 21014 19668 21020
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19260 20466 19288 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19444 19854 19472 20198
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19352 19378 19380 19722
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19168 18958 19288 18986
rect 19352 18970 19380 19314
rect 19260 18902 19288 18958
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18800 16590 18828 17478
rect 19260 16998 19288 18838
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18290 20024 21422
rect 20272 21078 20300 22066
rect 20260 21072 20312 21078
rect 20260 21014 20312 21020
rect 20364 20942 20392 22646
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20456 21010 20484 22510
rect 20548 21554 20576 23666
rect 20732 22778 20760 23802
rect 20916 23322 20944 24346
rect 21008 23798 21036 25842
rect 21744 25430 21772 26182
rect 22112 25922 22140 26454
rect 22204 26314 22232 26726
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22112 25894 22232 25922
rect 21732 25424 21784 25430
rect 21732 25366 21784 25372
rect 22204 24834 22232 25894
rect 22066 24818 22232 24834
rect 22054 24812 22232 24818
rect 22106 24806 22232 24812
rect 22054 24754 22106 24760
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 22112 24410 22140 24618
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 21284 23662 21312 24074
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20916 21622 20944 23122
rect 21008 22574 21036 23462
rect 21284 23118 21312 23598
rect 21732 23180 21784 23186
rect 21732 23122 21784 23128
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21284 22710 21312 23054
rect 21272 22704 21324 22710
rect 21272 22646 21324 22652
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20180 20262 20208 20878
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 20058 20392 20198
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19064 16720 19116 16726
rect 19064 16662 19116 16668
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 19076 16250 19104 16662
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18524 15609 18552 16118
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18800 15706 18828 16050
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18510 15600 18566 15609
rect 18510 15535 18566 15544
rect 19628 15502 19656 15982
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18248 14482 18276 14826
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 20088 14414 20116 19926
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20168 19440 20220 19446
rect 20272 19417 20300 19450
rect 20168 19382 20220 19388
rect 20258 19408 20314 19417
rect 20180 18766 20208 19382
rect 20258 19343 20314 19352
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18766 20392 19110
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18358 20300 18566
rect 20456 18426 20484 20946
rect 20548 20466 20576 21490
rect 21008 21146 21036 22510
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21560 22030 21588 22374
rect 21652 22234 21680 22578
rect 21744 22574 21772 23122
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21744 22030 21772 22510
rect 21836 22030 21864 22646
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21744 21622 21772 21966
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20916 20398 20944 20878
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20548 19174 20576 19858
rect 21008 19854 21036 20402
rect 21100 20058 21128 20878
rect 21284 20330 21312 21082
rect 21744 21010 21772 21558
rect 21836 21554 21864 21966
rect 22020 21690 22048 23734
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22204 22574 22232 23122
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 22204 21486 22232 22510
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22192 21072 22244 21078
rect 22112 21020 22192 21026
rect 22112 21014 22244 21020
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 22112 20998 22232 21014
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21468 20602 21496 20742
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20640 19446 20668 19790
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20994 19408 21050 19417
rect 20994 19343 20996 19352
rect 21048 19343 21050 19352
rect 20996 19314 21048 19320
rect 21100 19310 21128 19994
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 21192 18766 21220 19790
rect 21284 19718 21312 20266
rect 21376 20058 21404 20402
rect 22112 20262 22140 20998
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 22112 19378 22140 20198
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 21376 18970 21404 19314
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 22020 18766 22048 19110
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20732 18426 20760 18634
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 22296 16182 22324 26794
rect 22388 24410 22416 27118
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 22480 25430 22508 25842
rect 22468 25424 22520 25430
rect 22572 25401 22600 30194
rect 23032 29646 23060 30738
rect 23124 30394 23152 31282
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 23112 30388 23164 30394
rect 23112 30330 23164 30336
rect 23020 29640 23072 29646
rect 23020 29582 23072 29588
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 22756 28082 22784 29174
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 22928 29096 22980 29102
rect 22928 29038 22980 29044
rect 22940 28694 22968 29038
rect 22928 28688 22980 28694
rect 22928 28630 22980 28636
rect 23020 28620 23072 28626
rect 23020 28562 23072 28568
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22664 27470 22692 27814
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22664 25702 22692 27406
rect 22756 25838 22784 28018
rect 22744 25832 22796 25838
rect 22744 25774 22796 25780
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22468 25366 22520 25372
rect 22558 25392 22614 25401
rect 22558 25327 22614 25336
rect 22664 24886 22692 25638
rect 23032 25498 23060 28562
rect 23124 28422 23152 29106
rect 23216 28558 23244 31078
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 23308 29782 23336 30126
rect 23400 29850 23428 31282
rect 24768 31272 24820 31278
rect 24768 31214 24820 31220
rect 24676 31136 24728 31142
rect 24676 31078 24728 31084
rect 24688 30938 24716 31078
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24688 30394 24716 30670
rect 24676 30388 24728 30394
rect 24676 30330 24728 30336
rect 24584 30184 24636 30190
rect 24584 30126 24636 30132
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23296 29776 23348 29782
rect 23296 29718 23348 29724
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 23124 26926 23152 28358
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 23308 26466 23336 29718
rect 24308 28552 24360 28558
rect 24308 28494 24360 28500
rect 24320 28082 24348 28494
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24308 28076 24360 28082
rect 24308 28018 24360 28024
rect 24032 27872 24084 27878
rect 24032 27814 24084 27820
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23492 26518 23520 27474
rect 24044 27470 24072 27814
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24228 27130 24256 28018
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24412 26994 24440 27950
rect 23848 26988 23900 26994
rect 23848 26930 23900 26936
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 23216 26438 23336 26466
rect 23480 26512 23532 26518
rect 23480 26454 23532 26460
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22848 24954 22876 25298
rect 22836 24948 22888 24954
rect 22836 24890 22888 24896
rect 22652 24880 22704 24886
rect 22652 24822 22704 24828
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22388 23610 22416 24346
rect 23216 23730 23244 26438
rect 23492 25906 23520 26454
rect 23860 26042 23888 26930
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 24412 25906 24440 26930
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 24400 25900 24452 25906
rect 24400 25842 24452 25848
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 23308 23730 23336 25774
rect 23756 25696 23808 25702
rect 23756 25638 23808 25644
rect 23388 24948 23440 24954
rect 23388 24890 23440 24896
rect 23400 24206 23428 24890
rect 23768 24274 23796 25638
rect 24596 24818 24624 30126
rect 24688 29510 24716 30330
rect 24676 29504 24728 29510
rect 24676 29446 24728 29452
rect 24780 26874 24808 31214
rect 24872 29850 24900 31282
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 25056 30190 25084 30670
rect 25332 30326 25360 31350
rect 32968 31210 32996 37198
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 32956 31204 33008 31210
rect 32956 31146 33008 31152
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 25320 30320 25372 30326
rect 25320 30262 25372 30268
rect 25044 30184 25096 30190
rect 25096 30132 25176 30138
rect 25044 30126 25176 30132
rect 25056 30110 25176 30126
rect 25044 30048 25096 30054
rect 25044 29990 25096 29996
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 25056 29646 25084 29990
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 25056 29306 25084 29582
rect 25148 29578 25176 30110
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 25044 29300 25096 29306
rect 25044 29242 25096 29248
rect 25044 29096 25096 29102
rect 25044 29038 25096 29044
rect 25056 28762 25084 29038
rect 25044 28756 25096 28762
rect 25044 28698 25096 28704
rect 24860 28008 24912 28014
rect 24860 27950 24912 27956
rect 24872 27402 24900 27950
rect 25148 27606 25176 29514
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 37844 27606 37872 37198
rect 39316 37126 39344 39200
rect 39304 37120 39356 37126
rect 39304 37062 39356 37068
rect 38292 32904 38344 32910
rect 38292 32846 38344 32852
rect 38304 32745 38332 32846
rect 38290 32736 38346 32745
rect 38290 32671 38346 32680
rect 25136 27600 25188 27606
rect 25136 27542 25188 27548
rect 37832 27600 37884 27606
rect 37832 27542 37884 27548
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 24872 26994 24900 27338
rect 24952 27056 25004 27062
rect 24952 26998 25004 27004
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24688 26846 24808 26874
rect 24688 25838 24716 26846
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 24780 26382 24808 26726
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24964 26042 24992 26998
rect 25056 26586 25084 27474
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 26858 38056 27406
rect 38016 26852 38068 26858
rect 38016 26794 38068 26800
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 37188 26376 37240 26382
rect 37740 26376 37792 26382
rect 37188 26318 37240 26324
rect 37738 26344 37740 26353
rect 37792 26344 37794 26353
rect 24952 26036 25004 26042
rect 24952 25978 25004 25984
rect 37200 25945 37228 26318
rect 37738 26279 37794 26288
rect 37186 25936 37242 25945
rect 37186 25871 37242 25880
rect 24676 25832 24728 25838
rect 24676 25774 24728 25780
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24584 24812 24636 24818
rect 24584 24754 24636 24760
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23400 23866 23428 24142
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 22388 23594 22508 23610
rect 22388 23588 22520 23594
rect 22388 23582 22468 23588
rect 22468 23530 22520 23536
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22388 23118 22416 23462
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 23216 22030 23244 23666
rect 23492 23594 23520 24074
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23492 22778 23520 23530
rect 23952 23322 23980 23666
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23216 21690 23244 21966
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23032 21146 23060 21490
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22940 20466 22968 20742
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22756 19854 22784 20198
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18616 12986 18644 14282
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 19352 2650 19380 12786
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19444 2514 19472 14214
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 24780 2514 24808 24822
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 38292 19168 38344 19174
rect 38290 19136 38292 19145
rect 38344 19136 38346 19145
rect 34934 19068 35242 19077
rect 38290 19071 38346 19080
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 38292 12844 38344 12850
rect 38292 12786 38344 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 38304 12345 38332 12786
rect 38290 12336 38346 12345
rect 38290 12271 38346 12280
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 37556 5704 37608 5710
rect 37556 5646 37608 5652
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 37568 2922 37596 5646
rect 38200 5568 38252 5574
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 38198 5471 38254 5480
rect 37556 2916 37608 2922
rect 37556 2858 37608 2864
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 25884 2446 25912 2790
rect 32324 2446 32352 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 32 800 60 2382
rect 6472 800 6500 2382
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 800 12940 2246
rect 19352 800 19380 2382
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 25792 800 25820 2246
rect 32232 800 32260 2246
rect 38672 800 38700 2246
rect 18 200 74 800
rect 6458 200 6514 800
rect 12898 200 12954 800
rect 19338 200 19394 800
rect 25778 200 25834 800
rect 32218 200 32274 800
rect 38658 200 38714 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1766 34040 1822 34096
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 1766 27276 1768 27296
rect 1768 27276 1820 27296
rect 1820 27276 1822 27296
rect 1766 27240 1822 27276
rect 1766 20440 1822 20496
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 2042 26988 2098 27024
rect 2042 26968 2044 26988
rect 2044 26968 2096 26988
rect 2096 26968 2098 26988
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 6734 20984 6790 21040
rect 9862 30776 9918 30832
rect 10966 29028 11022 29064
rect 10966 29008 10968 29028
rect 10968 29008 11020 29028
rect 11020 29008 11022 29028
rect 9862 26288 9918 26344
rect 10414 25064 10470 25120
rect 8758 20984 8814 21040
rect 8022 19216 8078 19272
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1766 13676 1768 13696
rect 1768 13676 1820 13696
rect 1820 13676 1822 13696
rect 1766 13640 1822 13676
rect 1766 6840 1822 6896
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 10414 19216 10470 19272
rect 11058 18536 11114 18592
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9954 15444 9956 15464
rect 9956 15444 10008 15464
rect 10008 15444 10010 15464
rect 9954 15408 10010 15444
rect 10598 15000 10654 15056
rect 11242 15564 11298 15600
rect 11702 26560 11758 26616
rect 13174 30776 13230 30832
rect 13450 27512 13506 27568
rect 11242 15544 11244 15564
rect 11244 15544 11296 15564
rect 11296 15544 11298 15564
rect 11794 15136 11850 15192
rect 11978 15444 11980 15464
rect 11980 15444 12032 15464
rect 12032 15444 12034 15464
rect 11978 15408 12034 15444
rect 14646 31764 14648 31784
rect 14648 31764 14700 31784
rect 14700 31764 14702 31784
rect 14646 31728 14702 31764
rect 14922 31864 14978 31920
rect 13726 26696 13782 26752
rect 14830 27412 14832 27432
rect 14832 27412 14884 27432
rect 14884 27412 14886 27432
rect 14830 27376 14886 27412
rect 14922 26968 14978 27024
rect 14646 26696 14702 26752
rect 14278 23860 14334 23896
rect 14278 23840 14280 23860
rect 14280 23840 14332 23860
rect 14332 23840 14334 23860
rect 14738 26288 14794 26344
rect 14278 20460 14334 20496
rect 14278 20440 14280 20460
rect 14280 20440 14332 20460
rect 14332 20440 14334 20460
rect 14462 20168 14518 20224
rect 14922 25100 14924 25120
rect 14924 25100 14976 25120
rect 14976 25100 14978 25120
rect 14922 25064 14978 25100
rect 14922 23704 14978 23760
rect 16210 33396 16212 33416
rect 16212 33396 16264 33416
rect 16264 33396 16266 33416
rect 16210 33360 16266 33396
rect 15842 31884 15898 31920
rect 15842 31864 15844 31884
rect 15844 31864 15896 31884
rect 15896 31864 15898 31884
rect 15474 26732 15476 26752
rect 15476 26732 15528 26752
rect 15528 26732 15530 26752
rect 15474 26696 15530 26732
rect 16486 29688 16542 29744
rect 16210 27548 16212 27568
rect 16212 27548 16264 27568
rect 16264 27548 16266 27568
rect 16210 27512 16266 27548
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 17958 29044 17960 29064
rect 17960 29044 18012 29064
rect 18012 29044 18014 29064
rect 17958 29008 18014 29044
rect 16026 26308 16082 26344
rect 16026 26288 16028 26308
rect 16028 26288 16080 26308
rect 16080 26288 16082 26308
rect 15382 24656 15438 24712
rect 15658 24112 15714 24168
rect 16210 24928 16266 24984
rect 16670 26560 16726 26616
rect 15014 20304 15070 20360
rect 15658 19508 15714 19544
rect 15658 19488 15660 19508
rect 15660 19488 15712 19508
rect 15712 19488 15714 19508
rect 16302 23568 16358 23624
rect 16302 19488 16358 19544
rect 15566 16652 15622 16688
rect 15566 16632 15568 16652
rect 15568 16632 15620 16652
rect 15620 16632 15622 16652
rect 14278 15136 14334 15192
rect 14554 15020 14610 15056
rect 14554 15000 14556 15020
rect 14556 15000 14608 15020
rect 14608 15000 14610 15020
rect 17130 26696 17186 26752
rect 17038 26560 17094 26616
rect 16762 23840 16818 23896
rect 16854 20440 16910 20496
rect 17130 18572 17132 18592
rect 17132 18572 17184 18592
rect 17184 18572 17186 18592
rect 17130 18536 17186 18572
rect 17590 23568 17646 23624
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 17774 20168 17830 20224
rect 18326 20168 18382 20224
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19338 25372 19340 25392
rect 19340 25372 19392 25392
rect 19392 25372 19394 25392
rect 19338 25336 19394 25372
rect 19706 25220 19762 25256
rect 19706 25200 19708 25220
rect 19708 25200 19760 25220
rect 19760 25200 19762 25220
rect 19338 25064 19394 25120
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19154 24656 19210 24712
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 18510 15544 18566 15600
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20258 19352 20314 19408
rect 20994 19372 21050 19408
rect 20994 19352 20996 19372
rect 20996 19352 21048 19372
rect 21048 19352 21050 19372
rect 22558 25336 22614 25392
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 38290 32680 38346 32736
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 37738 26324 37740 26344
rect 37740 26324 37792 26344
rect 37792 26324 37794 26344
rect 37738 26288 37794 26324
rect 37186 25880 37242 25936
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 38290 19116 38292 19136
rect 38292 19116 38344 19136
rect 38344 19116 38346 19136
rect 38290 19080 38346 19116
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 38290 12280 38346 12336
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 16205 33420 16271 33421
rect 16205 33418 16252 33420
rect 16160 33416 16252 33418
rect 16160 33360 16210 33416
rect 16160 33358 16252 33360
rect 16205 33356 16252 33358
rect 16316 33356 16322 33420
rect 16205 33355 16271 33356
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 38285 32738 38351 32741
rect 39200 32738 39800 32768
rect 38285 32736 39800 32738
rect 38285 32680 38290 32736
rect 38346 32680 39800 32736
rect 38285 32678 39800 32680
rect 38285 32675 38351 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 14917 31922 14983 31925
rect 15837 31922 15903 31925
rect 14917 31920 15903 31922
rect 14917 31864 14922 31920
rect 14978 31864 15842 31920
rect 15898 31864 15903 31920
rect 14917 31862 15903 31864
rect 14917 31859 14983 31862
rect 15837 31859 15903 31862
rect 14641 31786 14707 31789
rect 14774 31786 14780 31788
rect 14641 31784 14780 31786
rect 14641 31728 14646 31784
rect 14702 31728 14780 31784
rect 14641 31726 14780 31728
rect 14641 31723 14707 31726
rect 14774 31724 14780 31726
rect 14844 31724 14850 31788
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 9857 30834 9923 30837
rect 13169 30834 13235 30837
rect 9857 30832 13235 30834
rect 9857 30776 9862 30832
rect 9918 30776 13174 30832
rect 13230 30776 13235 30832
rect 9857 30774 13235 30776
rect 9857 30771 9923 30774
rect 13169 30771 13235 30774
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 16481 29748 16547 29749
rect 16430 29684 16436 29748
rect 16500 29746 16547 29748
rect 16500 29744 16592 29746
rect 16542 29688 16592 29744
rect 16500 29686 16592 29688
rect 16500 29684 16547 29686
rect 16481 29683 16547 29684
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 10961 29066 11027 29069
rect 17953 29066 18019 29069
rect 10961 29064 18019 29066
rect 10961 29008 10966 29064
rect 11022 29008 17958 29064
rect 18014 29008 18019 29064
rect 10961 29006 18019 29008
rect 10961 29003 11027 29006
rect 17953 29003 18019 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 13445 27570 13511 27573
rect 16205 27570 16271 27573
rect 13445 27568 16271 27570
rect 13445 27512 13450 27568
rect 13506 27512 16210 27568
rect 16266 27512 16271 27568
rect 13445 27510 16271 27512
rect 13445 27507 13511 27510
rect 16205 27507 16271 27510
rect 14825 27434 14891 27437
rect 14958 27434 14964 27436
rect 14825 27432 14964 27434
rect 14825 27376 14830 27432
rect 14886 27376 14964 27432
rect 14825 27374 14964 27376
rect 14825 27371 14891 27374
rect 14958 27372 14964 27374
rect 15028 27372 15034 27436
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 2037 27026 2103 27029
rect 14917 27026 14983 27029
rect 2037 27024 14983 27026
rect 2037 26968 2042 27024
rect 2098 26968 14922 27024
rect 14978 26968 14983 27024
rect 2037 26966 14983 26968
rect 2037 26963 2103 26966
rect 14917 26963 14983 26966
rect 13721 26754 13787 26757
rect 14641 26754 14707 26757
rect 15469 26754 15535 26757
rect 17125 26754 17191 26757
rect 13721 26752 17191 26754
rect 13721 26696 13726 26752
rect 13782 26696 14646 26752
rect 14702 26696 15474 26752
rect 15530 26696 17130 26752
rect 17186 26696 17191 26752
rect 13721 26694 17191 26696
rect 13721 26691 13787 26694
rect 14641 26691 14707 26694
rect 15469 26691 15535 26694
rect 17125 26691 17191 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 11697 26618 11763 26621
rect 16665 26618 16731 26621
rect 17033 26618 17099 26621
rect 11697 26616 17099 26618
rect 11697 26560 11702 26616
rect 11758 26560 16670 26616
rect 16726 26560 17038 26616
rect 17094 26560 17099 26616
rect 11697 26558 17099 26560
rect 11697 26555 11763 26558
rect 16665 26555 16731 26558
rect 17033 26555 17099 26558
rect 9857 26346 9923 26349
rect 14733 26346 14799 26349
rect 9857 26344 14799 26346
rect 9857 26288 9862 26344
rect 9918 26288 14738 26344
rect 14794 26288 14799 26344
rect 9857 26286 14799 26288
rect 9857 26283 9923 26286
rect 14733 26283 14799 26286
rect 16021 26346 16087 26349
rect 37733 26346 37799 26349
rect 16021 26344 37799 26346
rect 16021 26288 16026 26344
rect 16082 26288 37738 26344
rect 37794 26288 37799 26344
rect 16021 26286 37799 26288
rect 16021 26283 16087 26286
rect 37733 26283 37799 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 37181 25938 37247 25941
rect 39200 25938 39800 25968
rect 37181 25936 39800 25938
rect 37181 25880 37186 25936
rect 37242 25880 39800 25936
rect 37181 25878 39800 25880
rect 37181 25875 37247 25878
rect 39200 25848 39800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19333 25394 19399 25397
rect 22553 25394 22619 25397
rect 19333 25392 22619 25394
rect 19333 25336 19338 25392
rect 19394 25336 22558 25392
rect 22614 25336 22619 25392
rect 19333 25334 22619 25336
rect 19333 25331 19399 25334
rect 22553 25331 22619 25334
rect 19701 25258 19767 25261
rect 19382 25256 19767 25258
rect 19382 25200 19706 25256
rect 19762 25200 19767 25256
rect 19382 25198 19767 25200
rect 19382 25125 19442 25198
rect 19701 25195 19767 25198
rect 10409 25122 10475 25125
rect 14917 25122 14983 25125
rect 10409 25120 14983 25122
rect 10409 25064 10414 25120
rect 10470 25064 14922 25120
rect 14978 25064 14983 25120
rect 10409 25062 14983 25064
rect 10409 25059 10475 25062
rect 14917 25059 14983 25062
rect 19333 25120 19442 25125
rect 19333 25064 19338 25120
rect 19394 25064 19442 25120
rect 19333 25062 19442 25064
rect 19333 25059 19399 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 15694 24924 15700 24988
rect 15764 24986 15770 24988
rect 16205 24986 16271 24989
rect 15764 24984 16271 24986
rect 15764 24928 16210 24984
rect 16266 24928 16271 24984
rect 15764 24926 16271 24928
rect 15764 24924 15770 24926
rect 16205 24923 16271 24926
rect 15377 24714 15443 24717
rect 19149 24714 19215 24717
rect 15377 24712 19215 24714
rect 15377 24656 15382 24712
rect 15438 24656 19154 24712
rect 19210 24656 19215 24712
rect 15377 24654 19215 24656
rect 15377 24651 15443 24654
rect 19149 24651 19215 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 14774 24108 14780 24172
rect 14844 24170 14850 24172
rect 15653 24170 15719 24173
rect 14844 24168 15719 24170
rect 14844 24112 15658 24168
rect 15714 24112 15719 24168
rect 14844 24110 15719 24112
rect 14844 24108 14850 24110
rect 15653 24107 15719 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 14273 23898 14339 23901
rect 16430 23898 16436 23900
rect 14273 23896 16436 23898
rect 14273 23840 14278 23896
rect 14334 23840 16436 23896
rect 14273 23838 16436 23840
rect 14273 23835 14339 23838
rect 14920 23765 14980 23838
rect 16430 23836 16436 23838
rect 16500 23898 16506 23900
rect 16757 23898 16823 23901
rect 16500 23896 16823 23898
rect 16500 23840 16762 23896
rect 16818 23840 16823 23896
rect 16500 23838 16823 23840
rect 16500 23836 16506 23838
rect 16757 23835 16823 23838
rect 14917 23760 14983 23765
rect 14917 23704 14922 23760
rect 14978 23704 14983 23760
rect 14917 23699 14983 23704
rect 16297 23626 16363 23629
rect 17585 23626 17651 23629
rect 16297 23624 17651 23626
rect 16297 23568 16302 23624
rect 16358 23568 17590 23624
rect 17646 23568 17651 23624
rect 16297 23566 17651 23568
rect 16297 23563 16363 23566
rect 17585 23563 17651 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 6729 21042 6795 21045
rect 8753 21042 8819 21045
rect 6729 21040 8819 21042
rect 6729 20984 6734 21040
rect 6790 20984 8758 21040
rect 8814 20984 8819 21040
rect 6729 20982 8819 20984
rect 6729 20979 6795 20982
rect 8753 20979 8819 20982
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 14273 20498 14339 20501
rect 16849 20498 16915 20501
rect 14273 20496 16915 20498
rect 14273 20440 14278 20496
rect 14334 20440 16854 20496
rect 16910 20440 16915 20496
rect 14273 20438 16915 20440
rect 14273 20435 14339 20438
rect 16849 20435 16915 20438
rect 15009 20364 15075 20365
rect 14958 20362 14964 20364
rect 14918 20302 14964 20362
rect 15028 20360 15075 20364
rect 15070 20304 15075 20360
rect 14958 20300 14964 20302
rect 15028 20300 15075 20304
rect 15009 20299 15075 20300
rect 14457 20226 14523 20229
rect 17769 20226 17835 20229
rect 18321 20226 18387 20229
rect 14457 20224 18387 20226
rect 14457 20168 14462 20224
rect 14518 20168 17774 20224
rect 17830 20168 18326 20224
rect 18382 20168 18387 20224
rect 14457 20166 18387 20168
rect 14457 20163 14523 20166
rect 17769 20163 17835 20166
rect 18321 20163 18387 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 15653 19546 15719 19549
rect 16297 19546 16363 19549
rect 15653 19544 16363 19546
rect 15653 19488 15658 19544
rect 15714 19488 16302 19544
rect 16358 19488 16363 19544
rect 15653 19486 16363 19488
rect 15653 19483 15719 19486
rect 16297 19483 16363 19486
rect 20253 19410 20319 19413
rect 20989 19410 21055 19413
rect 20253 19408 21055 19410
rect 20253 19352 20258 19408
rect 20314 19352 20994 19408
rect 21050 19352 21055 19408
rect 20253 19350 21055 19352
rect 20253 19347 20319 19350
rect 20989 19347 21055 19350
rect 8017 19274 8083 19277
rect 10409 19274 10475 19277
rect 8017 19272 10475 19274
rect 8017 19216 8022 19272
rect 8078 19216 10414 19272
rect 10470 19216 10475 19272
rect 8017 19214 10475 19216
rect 8017 19211 8083 19214
rect 10409 19211 10475 19214
rect 38285 19138 38351 19141
rect 39200 19138 39800 19168
rect 38285 19136 39800 19138
rect 38285 19080 38290 19136
rect 38346 19080 39800 19136
rect 38285 19078 39800 19080
rect 38285 19075 38351 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 11053 18594 11119 18597
rect 16246 18594 16252 18596
rect 11053 18592 16252 18594
rect 11053 18536 11058 18592
rect 11114 18536 16252 18592
rect 11053 18534 16252 18536
rect 11053 18531 11119 18534
rect 16246 18532 16252 18534
rect 16316 18594 16322 18596
rect 17125 18594 17191 18597
rect 16316 18592 17191 18594
rect 16316 18536 17130 18592
rect 17186 18536 17191 18592
rect 16316 18534 17191 18536
rect 16316 18532 16322 18534
rect 17125 18531 17191 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 15561 16690 15627 16693
rect 15694 16690 15700 16692
rect 15561 16688 15700 16690
rect 15561 16632 15566 16688
rect 15622 16632 15700 16688
rect 15561 16630 15700 16632
rect 15561 16627 15627 16630
rect 15694 16628 15700 16630
rect 15764 16628 15770 16692
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 11237 15602 11303 15605
rect 18505 15602 18571 15605
rect 11237 15600 18571 15602
rect 11237 15544 11242 15600
rect 11298 15544 18510 15600
rect 18566 15544 18571 15600
rect 11237 15542 18571 15544
rect 11237 15539 11303 15542
rect 18505 15539 18571 15542
rect 9949 15466 10015 15469
rect 11973 15466 12039 15469
rect 9949 15464 12039 15466
rect 9949 15408 9954 15464
rect 10010 15408 11978 15464
rect 12034 15408 12039 15464
rect 9949 15406 12039 15408
rect 9949 15403 10015 15406
rect 11973 15403 12039 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 11789 15194 11855 15197
rect 14273 15194 14339 15197
rect 11789 15192 14339 15194
rect 11789 15136 11794 15192
rect 11850 15136 14278 15192
rect 14334 15136 14339 15192
rect 11789 15134 14339 15136
rect 11789 15131 11855 15134
rect 14273 15131 14339 15134
rect 10593 15058 10659 15061
rect 14549 15058 14615 15061
rect 10593 15056 14615 15058
rect 10593 15000 10598 15056
rect 10654 15000 14554 15056
rect 14610 15000 14615 15056
rect 10593 14998 14615 15000
rect 10593 14995 10659 14998
rect 14549 14995 14615 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 38285 12338 38351 12341
rect 39200 12338 39800 12368
rect 38285 12336 39800 12338
rect 38285 12280 38290 12336
rect 38346 12280 39800 12336
rect 38285 12278 39800 12280
rect 38285 12275 38351 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1761 6898 1827 6901
rect 200 6896 1827 6898
rect 200 6840 1766 6896
rect 1822 6840 1827 6896
rect 200 6838 1827 6840
rect 200 6808 800 6838
rect 1761 6835 1827 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 16252 33416 16316 33420
rect 16252 33360 16266 33416
rect 16266 33360 16316 33416
rect 16252 33356 16316 33360
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 14780 31724 14844 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 16436 29744 16500 29748
rect 16436 29688 16486 29744
rect 16486 29688 16500 29744
rect 16436 29684 16500 29688
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 14964 27372 15028 27436
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 15700 24924 15764 24988
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 14780 24108 14844 24172
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 16436 23836 16500 23900
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 14964 20360 15028 20364
rect 14964 20304 15014 20360
rect 15014 20304 15028 20360
rect 14964 20300 15028 20304
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 16252 18532 16316 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 15700 16628 15764 16692
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 16251 33420 16317 33421
rect 16251 33356 16252 33420
rect 16316 33356 16317 33420
rect 16251 33355 16317 33356
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 14779 31788 14845 31789
rect 14779 31724 14780 31788
rect 14844 31724 14845 31788
rect 14779 31723 14845 31724
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 14782 24173 14842 31723
rect 14963 27436 15029 27437
rect 14963 27372 14964 27436
rect 15028 27372 15029 27436
rect 14963 27371 15029 27372
rect 14779 24172 14845 24173
rect 14779 24108 14780 24172
rect 14844 24108 14845 24172
rect 14779 24107 14845 24108
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 14966 20365 15026 27371
rect 15699 24988 15765 24989
rect 15699 24924 15700 24988
rect 15764 24924 15765 24988
rect 15699 24923 15765 24924
rect 14963 20364 15029 20365
rect 14963 20300 14964 20364
rect 15028 20300 15029 20364
rect 14963 20299 15029 20300
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 15702 16693 15762 24923
rect 16254 18597 16314 33355
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 16435 29748 16501 29749
rect 16435 29684 16436 29748
rect 16500 29684 16501 29748
rect 16435 29683 16501 29684
rect 16438 23901 16498 29683
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 16435 23900 16501 23901
rect 16435 23836 16436 23900
rect 16500 23836 16501 23900
rect 16435 23835 16501 23836
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 16251 18596 16317 18597
rect 16251 18532 16252 18596
rect 16316 18532 16317 18596
rect 16251 18531 16317 18532
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 15699 16692 15765 16693
rect 15699 16628 15700 16692
rect 15764 16628 15765 16692
rect 15699 16627 15765 16628
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32752 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform -1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1667941163
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1667941163
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1667941163
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1667941163
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1667941163
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1667941163
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1667941163
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1667941163
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1667941163
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1667941163
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_342
timestamp 1667941163
transform 1 0 32568 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_346
timestamp 1667941163
transform 1 0 32936 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_358
timestamp 1667941163
transform 1 0 34040 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_370
timestamp 1667941163
transform 1 0 35144 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1667941163
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_393
timestamp 1667941163
transform 1 0 37260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_397
timestamp 1667941163
transform 1 0 37628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_10
timestamp 1667941163
transform 1 0 2024 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1667941163
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_179
timestamp 1667941163
transform 1 0 17572 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_98
timestamp 1667941163
transform 1 0 10120 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_104
timestamp 1667941163
transform 1 0 10672 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1667941163
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1667941163
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1667941163
transform 1 0 14260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1667941163
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_158
timestamp 1667941163
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_192
timestamp 1667941163
transform 1 0 18768 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_204
timestamp 1667941163
transform 1 0 19872 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1667941163
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_107
timestamp 1667941163
transform 1 0 10948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_113
timestamp 1667941163
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1667941163
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1667941163
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_157
timestamp 1667941163
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_174
timestamp 1667941163
transform 1 0 17112 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1667941163
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_89
timestamp 1667941163
transform 1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1667941163
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_127
timestamp 1667941163
transform 1 0 12788 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_145
timestamp 1667941163
transform 1 0 14444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1667941163
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_158
timestamp 1667941163
transform 1 0 15640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1667941163
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_190
timestamp 1667941163
transform 1 0 18584 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_90
timestamp 1667941163
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_102
timestamp 1667941163
transform 1 0 10488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1667941163
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1667941163
transform 1 0 12328 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1667941163
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 1667941163
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_161
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_167
timestamp 1667941163
transform 1 0 16468 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_214
timestamp 1667941163
transform 1 0 20792 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_226
timestamp 1667941163
transform 1 0 21896 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_238
timestamp 1667941163
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1667941163
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1667941163
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_123
timestamp 1667941163
transform 1 0 12420 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_134
timestamp 1667941163
transform 1 0 13432 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_147
timestamp 1667941163
transform 1 0 14628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_158
timestamp 1667941163
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_176
timestamp 1667941163
transform 1 0 17296 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_190
timestamp 1667941163
transform 1 0 18584 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_202
timestamp 1667941163
transform 1 0 19688 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1667941163
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1667941163
transform 1 0 9660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_118
timestamp 1667941163
transform 1 0 11960 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_132
timestamp 1667941163
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_157
timestamp 1667941163
transform 1 0 15548 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_163
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_173
timestamp 1667941163
transform 1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1667941163
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_202
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_214
timestamp 1667941163
transform 1 0 20792 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_226
timestamp 1667941163
transform 1 0 21896 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_238
timestamp 1667941163
transform 1 0 23000 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_65
timestamp 1667941163
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_85
timestamp 1667941163
transform 1 0 8924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_90
timestamp 1667941163
transform 1 0 9384 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_102
timestamp 1667941163
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_122
timestamp 1667941163
transform 1 0 12328 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_131
timestamp 1667941163
transform 1 0 13156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_140
timestamp 1667941163
transform 1 0 13984 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1667941163
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_156
timestamp 1667941163
transform 1 0 15456 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1667941163
transform 1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_190
timestamp 1667941163
transform 1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_197
timestamp 1667941163
transform 1 0 19228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_209
timestamp 1667941163
transform 1 0 20332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1667941163
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_35
timestamp 1667941163
transform 1 0 4324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_47
timestamp 1667941163
transform 1 0 5428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_55
timestamp 1667941163
transform 1 0 6164 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_60
timestamp 1667941163
transform 1 0 6624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1667941163
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_103
timestamp 1667941163
transform 1 0 10580 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1667941163
transform 1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1667941163
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1667941163
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_162
timestamp 1667941163
transform 1 0 16008 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_169
timestamp 1667941163
transform 1 0 16652 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1667941163
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1667941163
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1667941163
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1667941163
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1667941163
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1667941163
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1667941163
transform 1 0 7544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_76
timestamp 1667941163
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_84
timestamp 1667941163
transform 1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_92
timestamp 1667941163
transform 1 0 9568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_99
timestamp 1667941163
transform 1 0 10212 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1667941163
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_139
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_158
timestamp 1667941163
transform 1 0 15640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1667941163
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_21
timestamp 1667941163
transform 1 0 3036 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 1667941163
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_47
timestamp 1667941163
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_51
timestamp 1667941163
transform 1 0 5796 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_59
timestamp 1667941163
transform 1 0 6532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_73
timestamp 1667941163
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1667941163
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_102
timestamp 1667941163
transform 1 0 10488 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_115
timestamp 1667941163
transform 1 0 11684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_126
timestamp 1667941163
transform 1 0 12696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1667941163
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1667941163
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_167
timestamp 1667941163
transform 1 0 16468 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1667941163
transform 1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_184
timestamp 1667941163
transform 1 0 18032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1667941163
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1667941163
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_24
timestamp 1667941163
transform 1 0 3312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_43
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_64
timestamp 1667941163
transform 1 0 6992 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_70
timestamp 1667941163
transform 1 0 7544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_78
timestamp 1667941163
transform 1 0 8280 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_82
timestamp 1667941163
transform 1 0 8648 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_99
timestamp 1667941163
transform 1 0 10212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1667941163
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1667941163
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_142
timestamp 1667941163
transform 1 0 14168 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_150
timestamp 1667941163
transform 1 0 14904 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_177
timestamp 1667941163
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_182
timestamp 1667941163
transform 1 0 17848 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_190
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1667941163
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1667941163
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_40
timestamp 1667941163
transform 1 0 4784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1667941163
transform 1 0 5888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1667941163
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_101
timestamp 1667941163
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_127
timestamp 1667941163
transform 1 0 12788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_131
timestamp 1667941163
transform 1 0 13156 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1667941163
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_149
timestamp 1667941163
transform 1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_157
timestamp 1667941163
transform 1 0 15548 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_163
timestamp 1667941163
transform 1 0 16100 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1667941163
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1667941163
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_186
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1667941163
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1667941163
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_210
timestamp 1667941163
transform 1 0 20424 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_234
timestamp 1667941163
transform 1 0 22632 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_17
timestamp 1667941163
transform 1 0 2668 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1667941163
transform 1 0 4784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp 1667941163
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_64
timestamp 1667941163
transform 1 0 6992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_68
timestamp 1667941163
transform 1 0 7360 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1667941163
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1667941163
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_104
timestamp 1667941163
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1667941163
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1667941163
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_139
timestamp 1667941163
transform 1 0 13892 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 1667941163
transform 1 0 14628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_155
timestamp 1667941163
transform 1 0 15364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_174
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1667941163
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_190
timestamp 1667941163
transform 1 0 18584 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1667941163
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_204
timestamp 1667941163
transform 1 0 19872 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_208
timestamp 1667941163
transform 1 0 20240 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_214
timestamp 1667941163
transform 1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_242
timestamp 1667941163
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1667941163
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_266
timestamp 1667941163
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_401
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1667941163
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_39
timestamp 1667941163
transform 1 0 4692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_51
timestamp 1667941163
transform 1 0 5796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1667941163
transform 1 0 6900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_70
timestamp 1667941163
transform 1 0 7544 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1667941163
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1667941163
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1667941163
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1667941163
transform 1 0 12972 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1667941163
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1667941163
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_171
timestamp 1667941163
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1667941163
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_207
timestamp 1667941163
transform 1 0 20148 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_220
timestamp 1667941163
transform 1 0 21344 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_226
timestamp 1667941163
transform 1 0 21896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1667941163
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_14
timestamp 1667941163
transform 1 0 2392 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_26
timestamp 1667941163
transform 1 0 3496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_36
timestamp 1667941163
transform 1 0 4416 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_44
timestamp 1667941163
transform 1 0 5152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_71
timestamp 1667941163
transform 1 0 7636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_83
timestamp 1667941163
transform 1 0 8740 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_96
timestamp 1667941163
transform 1 0 9936 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_122
timestamp 1667941163
transform 1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_133
timestamp 1667941163
transform 1 0 13340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_141
timestamp 1667941163
transform 1 0 14076 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_150
timestamp 1667941163
transform 1 0 14904 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_177
timestamp 1667941163
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_188
timestamp 1667941163
transform 1 0 18400 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1667941163
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1667941163
transform 1 0 20424 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1667941163
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_231
timestamp 1667941163
transform 1 0 22356 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_238
timestamp 1667941163
transform 1 0 23000 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_250
timestamp 1667941163
transform 1 0 24104 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_262
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1667941163
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_9
timestamp 1667941163
transform 1 0 1932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_16
timestamp 1667941163
transform 1 0 2576 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_22
timestamp 1667941163
transform 1 0 3128 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_39
timestamp 1667941163
transform 1 0 4692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_47
timestamp 1667941163
transform 1 0 5428 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_55
timestamp 1667941163
transform 1 0 6164 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_66
timestamp 1667941163
transform 1 0 7176 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1667941163
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_94
timestamp 1667941163
transform 1 0 9752 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_100
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp 1667941163
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1667941163
transform 1 0 11960 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_125
timestamp 1667941163
transform 1 0 12604 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_131
timestamp 1667941163
transform 1 0 13156 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1667941163
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1667941163
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_170
timestamp 1667941163
transform 1 0 16744 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_178
timestamp 1667941163
transform 1 0 17480 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1667941163
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_188
timestamp 1667941163
transform 1 0 18400 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1667941163
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_204
timestamp 1667941163
transform 1 0 19872 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_216
timestamp 1667941163
transform 1 0 20976 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_224
timestamp 1667941163
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1667941163
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1667941163
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_11
timestamp 1667941163
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_19
timestamp 1667941163
transform 1 0 2852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_30
timestamp 1667941163
transform 1 0 3864 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_34
timestamp 1667941163
transform 1 0 4232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_42
timestamp 1667941163
transform 1 0 4968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_46
timestamp 1667941163
transform 1 0 5336 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_63
timestamp 1667941163
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_67
timestamp 1667941163
transform 1 0 7268 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1667941163
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1667941163
transform 1 0 9016 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_95
timestamp 1667941163
transform 1 0 9844 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_103
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_126
timestamp 1667941163
transform 1 0 12696 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_138
timestamp 1667941163
transform 1 0 13800 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1667941163
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1667941163
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_190
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_198
timestamp 1667941163
transform 1 0 19320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_204
timestamp 1667941163
transform 1 0 19872 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_212
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1667941163
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1667941163
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_248
timestamp 1667941163
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_260
timestamp 1667941163
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1667941163
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_14
timestamp 1667941163
transform 1 0 2392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 1667941163
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_37
timestamp 1667941163
transform 1 0 4508 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_57
timestamp 1667941163
transform 1 0 6348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_69
timestamp 1667941163
transform 1 0 7452 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1667941163
transform 1 0 9476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_99
timestamp 1667941163
transform 1 0 10212 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_107
timestamp 1667941163
transform 1 0 10948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_116
timestamp 1667941163
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1667941163
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_159
timestamp 1667941163
transform 1 0 15732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_167
timestamp 1667941163
transform 1 0 16468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_185
timestamp 1667941163
transform 1 0 18124 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1667941163
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_219
timestamp 1667941163
transform 1 0 21252 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_226
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_230
timestamp 1667941163
transform 1 0 22264 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_241
timestamp 1667941163
transform 1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1667941163
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1667941163
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_29
timestamp 1667941163
transform 1 0 3772 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_36
timestamp 1667941163
transform 1 0 4416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_44
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_49
timestamp 1667941163
transform 1 0 5612 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_75
timestamp 1667941163
transform 1 0 8004 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_87
timestamp 1667941163
transform 1 0 9108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1667941163
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1667941163
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_133
timestamp 1667941163
transform 1 0 13340 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_138
timestamp 1667941163
transform 1 0 13800 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_150
timestamp 1667941163
transform 1 0 14904 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_173
timestamp 1667941163
transform 1 0 17020 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_182
timestamp 1667941163
transform 1 0 17848 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_194
timestamp 1667941163
transform 1 0 18952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_202
timestamp 1667941163
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_212
timestamp 1667941163
transform 1 0 20608 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_245
timestamp 1667941163
transform 1 0 23644 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_257
timestamp 1667941163
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1667941163
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1667941163
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_37
timestamp 1667941163
transform 1 0 4508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_45
timestamp 1667941163
transform 1 0 5244 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_51
timestamp 1667941163
transform 1 0 5796 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_55
timestamp 1667941163
transform 1 0 6164 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_63
timestamp 1667941163
transform 1 0 6900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_75
timestamp 1667941163
transform 1 0 8004 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_93
timestamp 1667941163
transform 1 0 9660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_105
timestamp 1667941163
transform 1 0 10764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_117
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_125
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_131
timestamp 1667941163
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_172
timestamp 1667941163
transform 1 0 16928 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_206
timestamp 1667941163
transform 1 0 20056 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_214
timestamp 1667941163
transform 1 0 20792 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_222
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1667941163
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1667941163
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_18
timestamp 1667941163
transform 1 0 2760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_29
timestamp 1667941163
transform 1 0 3772 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_47
timestamp 1667941163
transform 1 0 5428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_64
timestamp 1667941163
transform 1 0 6992 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_75
timestamp 1667941163
transform 1 0 8004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_95
timestamp 1667941163
transform 1 0 9844 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_127
timestamp 1667941163
transform 1 0 12788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_134
timestamp 1667941163
transform 1 0 13432 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_138
timestamp 1667941163
transform 1 0 13800 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_153
timestamp 1667941163
transform 1 0 15180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1667941163
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_201
timestamp 1667941163
transform 1 0 19596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_209
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_232
timestamp 1667941163
transform 1 0 22448 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_245
timestamp 1667941163
transform 1 0 23644 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_257
timestamp 1667941163
transform 1 0 24748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1667941163
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_39
timestamp 1667941163
transform 1 0 4692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_47
timestamp 1667941163
transform 1 0 5428 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_57
timestamp 1667941163
transform 1 0 6348 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1667941163
transform 1 0 7544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1667941163
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1667941163
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_110
timestamp 1667941163
transform 1 0 11224 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1667941163
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_131
timestamp 1667941163
transform 1 0 13156 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_159
timestamp 1667941163
transform 1 0 15732 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_169
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1667941163
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_207
timestamp 1667941163
transform 1 0 20148 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_218
timestamp 1667941163
transform 1 0 21160 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_227
timestamp 1667941163
transform 1 0 21988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_235
timestamp 1667941163
transform 1 0 22724 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1667941163
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1667941163
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_11
timestamp 1667941163
transform 1 0 2116 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_21
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_28
timestamp 1667941163
transform 1 0 3680 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_36
timestamp 1667941163
transform 1 0 4416 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1667941163
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_91
timestamp 1667941163
transform 1 0 9476 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1667941163
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_118
timestamp 1667941163
transform 1 0 11960 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_130
timestamp 1667941163
transform 1 0 13064 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1667941163
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_143
timestamp 1667941163
transform 1 0 14260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_183
timestamp 1667941163
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1667941163
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_206
timestamp 1667941163
transform 1 0 20056 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1667941163
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1667941163
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_244
timestamp 1667941163
transform 1 0 23552 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_252
timestamp 1667941163
transform 1 0 24288 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_258
timestamp 1667941163
transform 1 0 24840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1667941163
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_57
timestamp 1667941163
transform 1 0 6348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_63
timestamp 1667941163
transform 1 0 6900 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_73
timestamp 1667941163
transform 1 0 7820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_90
timestamp 1667941163
transform 1 0 9384 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1667941163
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_108
timestamp 1667941163
transform 1 0 11040 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_120
timestamp 1667941163
transform 1 0 12144 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_128
timestamp 1667941163
transform 1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1667941163
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_154
timestamp 1667941163
transform 1 0 15272 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_171
timestamp 1667941163
transform 1 0 16836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_181
timestamp 1667941163
transform 1 0 17756 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_202
timestamp 1667941163
transform 1 0 19688 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_208
timestamp 1667941163
transform 1 0 20240 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1667941163
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_240
timestamp 1667941163
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_18
timestamp 1667941163
transform 1 0 2760 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_35
timestamp 1667941163
transform 1 0 4324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_44
timestamp 1667941163
transform 1 0 5152 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1667941163
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_63
timestamp 1667941163
transform 1 0 6900 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_74
timestamp 1667941163
transform 1 0 7912 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_87
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_95
timestamp 1667941163
transform 1 0 9844 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1667941163
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_122
timestamp 1667941163
transform 1 0 12328 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_130
timestamp 1667941163
transform 1 0 13064 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_141
timestamp 1667941163
transform 1 0 14076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1667941163
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_154
timestamp 1667941163
transform 1 0 15272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1667941163
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_179
timestamp 1667941163
transform 1 0 17572 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_189
timestamp 1667941163
transform 1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1667941163
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_209
timestamp 1667941163
transform 1 0 20332 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1667941163
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_231
timestamp 1667941163
transform 1 0 22356 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_236
timestamp 1667941163
transform 1 0 22816 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_250
timestamp 1667941163
transform 1 0 24104 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_260
timestamp 1667941163
transform 1 0 25024 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_272
timestamp 1667941163
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1667941163
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_39
timestamp 1667941163
transform 1 0 4692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_49
timestamp 1667941163
transform 1 0 5612 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_63
timestamp 1667941163
transform 1 0 6900 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_67
timestamp 1667941163
transform 1 0 7268 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_76
timestamp 1667941163
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_107
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_122
timestamp 1667941163
transform 1 0 12328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_131
timestamp 1667941163
transform 1 0 13156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_151
timestamp 1667941163
transform 1 0 14996 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_158
timestamp 1667941163
transform 1 0 15640 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_167
timestamp 1667941163
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1667941163
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1667941163
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_204
timestamp 1667941163
transform 1 0 19872 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_212
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1667941163
transform 1 0 21988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_244
timestamp 1667941163
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_262
timestamp 1667941163
transform 1 0 25208 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_274
timestamp 1667941163
transform 1 0 26312 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_286
timestamp 1667941163
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_298
timestamp 1667941163
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_7
timestamp 1667941163
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_11
timestamp 1667941163
transform 1 0 2116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_23
timestamp 1667941163
transform 1 0 3220 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_28
timestamp 1667941163
transform 1 0 3680 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_37
timestamp 1667941163
transform 1 0 4508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_47
timestamp 1667941163
transform 1 0 5428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_75
timestamp 1667941163
transform 1 0 8004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_89
timestamp 1667941163
transform 1 0 9292 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_117
timestamp 1667941163
transform 1 0 11868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1667941163
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_132
timestamp 1667941163
transform 1 0 13248 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_139
timestamp 1667941163
transform 1 0 13892 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1667941163
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_157
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_175
timestamp 1667941163
transform 1 0 17204 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1667941163
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1667941163
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_218
timestamp 1667941163
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_231
timestamp 1667941163
transform 1 0 22356 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_243
timestamp 1667941163
transform 1 0 23460 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_256
timestamp 1667941163
transform 1 0 24656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_268
timestamp 1667941163
transform 1 0 25760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_18
timestamp 1667941163
transform 1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1667941163
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_51
timestamp 1667941163
transform 1 0 5796 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_63
timestamp 1667941163
transform 1 0 6900 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_74
timestamp 1667941163
transform 1 0 7912 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_92
timestamp 1667941163
transform 1 0 9568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_104
timestamp 1667941163
transform 1 0 10672 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_110
timestamp 1667941163
transform 1 0 11224 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_117
timestamp 1667941163
transform 1 0 11868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_125
timestamp 1667941163
transform 1 0 12604 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1667941163
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_164
timestamp 1667941163
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_168
timestamp 1667941163
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1667941163
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_203
timestamp 1667941163
transform 1 0 19780 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_214
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_220
timestamp 1667941163
transform 1 0 21344 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_228
timestamp 1667941163
transform 1 0 22080 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_240
timestamp 1667941163
transform 1 0 23184 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_262
timestamp 1667941163
transform 1 0 25208 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_274
timestamp 1667941163
transform 1 0 26312 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_286
timestamp 1667941163
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_298
timestamp 1667941163
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1667941163
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_397
timestamp 1667941163
transform 1 0 37628 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_402
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1667941163
transform 1 0 38456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_34
timestamp 1667941163
transform 1 0 4232 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_46
timestamp 1667941163
transform 1 0 5336 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1667941163
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_76
timestamp 1667941163
transform 1 0 8096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_83
timestamp 1667941163
transform 1 0 8740 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1667941163
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_100
timestamp 1667941163
transform 1 0 10304 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_122
timestamp 1667941163
transform 1 0 12328 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_130
timestamp 1667941163
transform 1 0 13064 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_148
timestamp 1667941163
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1667941163
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_177
timestamp 1667941163
transform 1 0 17388 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_184
timestamp 1667941163
transform 1 0 18032 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_188
timestamp 1667941163
transform 1 0 18400 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_195
timestamp 1667941163
transform 1 0 19044 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_199
timestamp 1667941163
transform 1 0 19412 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_204
timestamp 1667941163
transform 1 0 19872 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_214
timestamp 1667941163
transform 1 0 20792 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1667941163
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_232
timestamp 1667941163
transform 1 0 22448 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_244
timestamp 1667941163
transform 1 0 23552 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_248
timestamp 1667941163
transform 1 0 23920 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_253
timestamp 1667941163
transform 1 0 24380 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_260
timestamp 1667941163
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1667941163
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_39
timestamp 1667941163
transform 1 0 4692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_43
timestamp 1667941163
transform 1 0 5060 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_50
timestamp 1667941163
transform 1 0 5704 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_58
timestamp 1667941163
transform 1 0 6440 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_62
timestamp 1667941163
transform 1 0 6808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_66
timestamp 1667941163
transform 1 0 7176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_93
timestamp 1667941163
transform 1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_101
timestamp 1667941163
transform 1 0 10396 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_119
timestamp 1667941163
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_131
timestamp 1667941163
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_149
timestamp 1667941163
transform 1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_158
timestamp 1667941163
transform 1 0 15640 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_167
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_179
timestamp 1667941163
transform 1 0 17572 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_184
timestamp 1667941163
transform 1 0 18032 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1667941163
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_206
timestamp 1667941163
transform 1 0 20056 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_214
timestamp 1667941163
transform 1 0 20792 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_222
timestamp 1667941163
transform 1 0 21528 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_226
timestamp 1667941163
transform 1 0 21896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1667941163
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_262
timestamp 1667941163
transform 1 0 25208 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_274
timestamp 1667941163
transform 1 0 26312 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_286
timestamp 1667941163
transform 1 0 27416 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_298
timestamp 1667941163
transform 1 0 28520 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1667941163
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_34
timestamp 1667941163
transform 1 0 4232 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_38
timestamp 1667941163
transform 1 0 4600 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_49
timestamp 1667941163
transform 1 0 5612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_66
timestamp 1667941163
transform 1 0 7176 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_74
timestamp 1667941163
transform 1 0 7912 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_82
timestamp 1667941163
transform 1 0 8648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_99
timestamp 1667941163
transform 1 0 10212 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_118
timestamp 1667941163
transform 1 0 11960 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_126
timestamp 1667941163
transform 1 0 12696 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_134
timestamp 1667941163
transform 1 0 13432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_139
timestamp 1667941163
transform 1 0 13892 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1667941163
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1667941163
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_173
timestamp 1667941163
transform 1 0 17020 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1667941163
transform 1 0 17480 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_188
timestamp 1667941163
transform 1 0 18400 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_197
timestamp 1667941163
transform 1 0 19228 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_212
timestamp 1667941163
transform 1 0 20608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1667941163
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_232
timestamp 1667941163
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_243
timestamp 1667941163
transform 1 0 23460 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_251
timestamp 1667941163
transform 1 0 24196 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_259
timestamp 1667941163
transform 1 0 24932 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_271
timestamp 1667941163
transform 1 0 26036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_19
timestamp 1667941163
transform 1 0 2852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1667941163
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_38
timestamp 1667941163
transform 1 0 4600 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_61
timestamp 1667941163
transform 1 0 6716 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_67
timestamp 1667941163
transform 1 0 7268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_75
timestamp 1667941163
transform 1 0 8004 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1667941163
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_92
timestamp 1667941163
transform 1 0 9568 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_108
timestamp 1667941163
transform 1 0 11040 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_116
timestamp 1667941163
transform 1 0 11776 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_125
timestamp 1667941163
transform 1 0 12604 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1667941163
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_148
timestamp 1667941163
transform 1 0 14720 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_158
timestamp 1667941163
transform 1 0 15640 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_168
timestamp 1667941163
transform 1 0 16560 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_180
timestamp 1667941163
transform 1 0 17664 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_212
timestamp 1667941163
transform 1 0 20608 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_229
timestamp 1667941163
transform 1 0 22172 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_238
timestamp 1667941163
transform 1 0 23000 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1667941163
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_261
timestamp 1667941163
transform 1 0 25116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_273
timestamp 1667941163
transform 1 0 26220 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_285
timestamp 1667941163
transform 1 0 27324 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_297
timestamp 1667941163
transform 1 0 28428 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1667941163
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_11
timestamp 1667941163
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_30
timestamp 1667941163
transform 1 0 3864 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_42
timestamp 1667941163
transform 1 0 4968 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1667941163
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_63
timestamp 1667941163
transform 1 0 6900 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_72
timestamp 1667941163
transform 1 0 7728 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_87
timestamp 1667941163
transform 1 0 9108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_94
timestamp 1667941163
transform 1 0 9752 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_103
timestamp 1667941163
transform 1 0 10580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_129
timestamp 1667941163
transform 1 0 12972 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_133
timestamp 1667941163
transform 1 0 13340 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_138
timestamp 1667941163
transform 1 0 13800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_157
timestamp 1667941163
transform 1 0 15548 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_188
timestamp 1667941163
transform 1 0 18400 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_192
timestamp 1667941163
transform 1 0 18768 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_196
timestamp 1667941163
transform 1 0 19136 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_204
timestamp 1667941163
transform 1 0 19872 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1667941163
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_233
timestamp 1667941163
transform 1 0 22540 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_239
timestamp 1667941163
transform 1 0 23092 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_247
timestamp 1667941163
transform 1 0 23828 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_255
timestamp 1667941163
transform 1 0 24564 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_264
timestamp 1667941163
transform 1 0 25392 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1667941163
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_11
timestamp 1667941163
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1667941163
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_35
timestamp 1667941163
transform 1 0 4324 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_42
timestamp 1667941163
transform 1 0 4968 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_50
timestamp 1667941163
transform 1 0 5704 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_55
timestamp 1667941163
transform 1 0 6164 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_63
timestamp 1667941163
transform 1 0 6900 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_69
timestamp 1667941163
transform 1 0 7452 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_94
timestamp 1667941163
transform 1 0 9752 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_104
timestamp 1667941163
transform 1 0 10672 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_108
timestamp 1667941163
transform 1 0 11040 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_118
timestamp 1667941163
transform 1 0 11960 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1667941163
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_150
timestamp 1667941163
transform 1 0 14904 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1667941163
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_168
timestamp 1667941163
transform 1 0 16560 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_176
timestamp 1667941163
transform 1 0 17296 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_185
timestamp 1667941163
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1667941163
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_204
timestamp 1667941163
transform 1 0 19872 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_211
timestamp 1667941163
transform 1 0 20516 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_225
timestamp 1667941163
transform 1 0 21804 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1667941163
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_261
timestamp 1667941163
transform 1 0 25116 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_273
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_285
timestamp 1667941163
transform 1 0 27324 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_297
timestamp 1667941163
transform 1 0 28428 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1667941163
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_25
timestamp 1667941163
transform 1 0 3404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1667941163
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_63
timestamp 1667941163
transform 1 0 6900 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_70
timestamp 1667941163
transform 1 0 7544 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_82
timestamp 1667941163
transform 1 0 8648 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_90
timestamp 1667941163
transform 1 0 9384 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_98
timestamp 1667941163
transform 1 0 10120 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_124
timestamp 1667941163
transform 1 0 12512 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_135
timestamp 1667941163
transform 1 0 13524 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_147
timestamp 1667941163
transform 1 0 14628 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_159
timestamp 1667941163
transform 1 0 15732 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1667941163
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_179
timestamp 1667941163
transform 1 0 17572 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_199
timestamp 1667941163
transform 1 0 19412 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1667941163
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_233
timestamp 1667941163
transform 1 0 22540 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_243
timestamp 1667941163
transform 1 0 23460 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_251
timestamp 1667941163
transform 1 0 24196 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_258
timestamp 1667941163
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1667941163
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1667941163
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_47
timestamp 1667941163
transform 1 0 5428 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_54
timestamp 1667941163
transform 1 0 6072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_68
timestamp 1667941163
transform 1 0 7360 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_76
timestamp 1667941163
transform 1 0 8096 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_89
timestamp 1667941163
transform 1 0 9292 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_96
timestamp 1667941163
transform 1 0 9936 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_107
timestamp 1667941163
transform 1 0 10948 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_119
timestamp 1667941163
transform 1 0 12052 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_132
timestamp 1667941163
transform 1 0 13248 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_150
timestamp 1667941163
transform 1 0 14904 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_161
timestamp 1667941163
transform 1 0 15916 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_185
timestamp 1667941163
transform 1 0 18124 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_193
timestamp 1667941163
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_206
timestamp 1667941163
transform 1 0 20056 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_218
timestamp 1667941163
transform 1 0 21160 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_230
timestamp 1667941163
transform 1 0 22264 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_242
timestamp 1667941163
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1667941163
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_75
timestamp 1667941163
transform 1 0 8004 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_82
timestamp 1667941163
transform 1 0 8648 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_95
timestamp 1667941163
transform 1 0 9844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_102
timestamp 1667941163
transform 1 0 10488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_109
timestamp 1667941163
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_122
timestamp 1667941163
transform 1 0 12328 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_129
timestamp 1667941163
transform 1 0 12972 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_133
timestamp 1667941163
transform 1 0 13340 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_138
timestamp 1667941163
transform 1 0 13800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_152
timestamp 1667941163
transform 1 0 15088 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_163
timestamp 1667941163
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_176
timestamp 1667941163
transform 1 0 17296 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_183
timestamp 1667941163
transform 1 0 17940 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_195
timestamp 1667941163
transform 1 0 19044 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_207
timestamp 1667941163
transform 1 0 20148 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1667941163
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_72
timestamp 1667941163
transform 1 0 7728 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_76
timestamp 1667941163
transform 1 0 8096 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_105
timestamp 1667941163
transform 1 0 10764 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_116
timestamp 1667941163
transform 1 0 11776 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 1667941163
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_145
timestamp 1667941163
transform 1 0 14444 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_150
timestamp 1667941163
transform 1 0 14904 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_158
timestamp 1667941163
transform 1 0 15640 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_178
timestamp 1667941163
transform 1 0 17480 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1667941163
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_85
timestamp 1667941163
transform 1 0 8924 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_91
timestamp 1667941163
transform 1 0 9476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1667941163
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_121
timestamp 1667941163
transform 1 0 12236 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_132
timestamp 1667941163
transform 1 0 13248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_156
timestamp 1667941163
transform 1 0 15456 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1667941163
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_96
timestamp 1667941163
transform 1 0 9936 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_108
timestamp 1667941163
transform 1 0 11040 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_120
timestamp 1667941163
transform 1 0 12144 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_125
timestamp 1667941163
transform 1 0 12604 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1667941163
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_148
timestamp 1667941163
transform 1 0 14720 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_160
timestamp 1667941163
transform 1 0 15824 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_164
timestamp 1667941163
transform 1 0 16192 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_176
timestamp 1667941163
transform 1 0 17296 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_188
timestamp 1667941163
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1667941163
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1667941163
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1667941163
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_202
timestamp 1667941163
transform 1 0 19688 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1667941163
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_8
timestamp 1667941163
transform 1 0 1840 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1667941163
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1667941163
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1667941163
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_159
timestamp 1667941163
transform 1 0 15732 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1667941163
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1667941163
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1667941163
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1667941163
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1667941163
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_345
timestamp 1667941163
transform 1 0 32844 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1667941163
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _0502_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17020 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0503_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18584 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0504_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0505_
timestamp 1667941163
transform 1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0506_
timestamp 1667941163
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0507_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0508_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _0509_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14812 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 16928 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0511_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17572 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0512_
timestamp 1667941163
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0513_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17020 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0515_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0516_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16928 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _0517_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17204 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0518_
timestamp 1667941163
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0519_
timestamp 1667941163
transform 1 0 23552 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0520_
timestamp 1667941163
transform 1 0 20884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0521_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0522_
timestamp 1667941163
transform 1 0 20608 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0523_
timestamp 1667941163
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _0524_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19688 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0525_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15272 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0526_
timestamp 1667941163
transform 1 0 15088 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0527_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14444 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0528_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0529_
timestamp 1667941163
transform 1 0 14260 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0530_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16008 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0531_
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0532_
timestamp 1667941163
transform 1 0 13248 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0533_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18308 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0534_
timestamp 1667941163
transform 1 0 15272 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0535_
timestamp 1667941163
transform 1 0 16928 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0536_
timestamp 1667941163
transform 1 0 14168 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0537_
timestamp 1667941163
transform 1 0 14168 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0538_
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0539_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15180 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0540_
timestamp 1667941163
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0541_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0542_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24380 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0543_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 15272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0545_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0546_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14444 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0547_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0548_
timestamp 1667941163
transform 1 0 13248 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0549_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0550_
timestamp 1667941163
transform 1 0 18492 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0551_
timestamp 1667941163
transform 1 0 19136 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0552_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0554_
timestamp 1667941163
transform 1 0 22448 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 23368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0556_
timestamp 1667941163
transform 1 0 24380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 21160 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 17756 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0559_
timestamp 1667941163
transform 1 0 20884 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0560_
timestamp 1667941163
transform 1 0 18492 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0561_
timestamp 1667941163
transform 1 0 18400 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0562_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0563_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20976 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0564_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20240 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0565_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0566_
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0567_
timestamp 1667941163
transform 1 0 23552 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0568_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0569_
timestamp 1667941163
transform 1 0 21988 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0570_
timestamp 1667941163
transform 1 0 22448 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0571_
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0572_
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0573_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0574_
timestamp 1667941163
transform 1 0 21988 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0575_
timestamp 1667941163
transform 1 0 24472 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0576_
timestamp 1667941163
transform 1 0 23644 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0577_
timestamp 1667941163
transform 1 0 17112 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0578_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0579_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0580_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0581_
timestamp 1667941163
transform 1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0582_
timestamp 1667941163
transform 1 0 22908 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0583_
timestamp 1667941163
transform 1 0 23184 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0584_
timestamp 1667941163
transform 1 0 24564 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0585_
timestamp 1667941163
transform 1 0 20148 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0586_
timestamp 1667941163
transform 1 0 20884 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0587_
timestamp 1667941163
transform 1 0 22816 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0588_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0589_
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0590_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0591_
timestamp 1667941163
transform 1 0 24288 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0592_
timestamp 1667941163
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0593_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24656 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0594_
timestamp 1667941163
transform 1 0 24380 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0595_
timestamp 1667941163
transform 1 0 6440 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0596_
timestamp 1667941163
transform 1 0 6624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0597_
timestamp 1667941163
transform 1 0 9108 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0598_
timestamp 1667941163
transform 1 0 10856 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0599_
timestamp 1667941163
transform 1 0 7268 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0600_
timestamp 1667941163
transform 1 0 3864 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0601_
timestamp 1667941163
transform 1 0 8096 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0602_
timestamp 1667941163
transform 1 0 7912 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0603_
timestamp 1667941163
transform 1 0 9108 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0604_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0605_
timestamp 1667941163
transform 1 0 4324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0606_
timestamp 1667941163
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0607_
timestamp 1667941163
transform 1 0 7912 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0608_
timestamp 1667941163
transform 1 0 7360 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0609_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7544 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0610_
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0611_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0612_
timestamp 1667941163
transform 1 0 23000 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0613_
timestamp 1667941163
transform 1 0 19412 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _0614_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15456 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_1  _0615_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17572 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0616_
timestamp 1667941163
transform 1 0 15456 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0617_
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0618_
timestamp 1667941163
transform 1 0 14168 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0619_
timestamp 1667941163
transform 1 0 14812 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0620_
timestamp 1667941163
transform 1 0 9936 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0621_
timestamp 1667941163
transform 1 0 15732 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0622_
timestamp 1667941163
transform 1 0 17940 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0623_
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0624_
timestamp 1667941163
transform 1 0 16008 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0625_
timestamp 1667941163
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0626_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0627_
timestamp 1667941163
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0628_
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0629_
timestamp 1667941163
transform 1 0 10304 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0630_
timestamp 1667941163
transform 1 0 18768 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0631_
timestamp 1667941163
transform 1 0 17388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0632_
timestamp 1667941163
transform 1 0 17848 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0633_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17848 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1667941163
transform 1 0 17848 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0635_
timestamp 1667941163
transform 1 0 19412 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0636_
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0637_
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1667941163
transform 1 0 19780 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1667941163
transform 1 0 20976 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0640_
timestamp 1667941163
transform 1 0 20056 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0641_
timestamp 1667941163
transform 1 0 19964 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 20240 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0643_
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0644_
timestamp 1667941163
transform 1 0 22080 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0645_
timestamp 1667941163
transform 1 0 10580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0646_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0647_
timestamp 1667941163
transform 1 0 16652 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0648_
timestamp 1667941163
transform 1 0 15824 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0649_
timestamp 1667941163
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0650_
timestamp 1667941163
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0652_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16560 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0653_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0654_
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0655_
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0656_
timestamp 1667941163
transform 1 0 18400 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0658_
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0659_
timestamp 1667941163
transform 1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0660_
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0661_
timestamp 1667941163
transform 1 0 10856 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0662_
timestamp 1667941163
transform 1 0 10856 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0663_
timestamp 1667941163
transform 1 0 9108 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0664_
timestamp 1667941163
transform 1 0 9936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0665_
timestamp 1667941163
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0666_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14352 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0667_
timestamp 1667941163
transform 1 0 10304 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0668_
timestamp 1667941163
transform 1 0 15088 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0669_
timestamp 1667941163
transform 1 0 14996 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 1667941163
transform 1 0 14628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0671_
timestamp 1667941163
transform 1 0 12328 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0673_
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0674_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0675_
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0677_
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0678_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10764 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0679_
timestamp 1667941163
transform 1 0 12696 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0680_
timestamp 1667941163
transform 1 0 11500 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0681_
timestamp 1667941163
transform 1 0 11316 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0682_
timestamp 1667941163
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0683_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11684 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0684_
timestamp 1667941163
transform 1 0 10580 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0685_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0686_
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0687_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0688_
timestamp 1667941163
transform 1 0 10304 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0689_
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0690_
timestamp 1667941163
transform 1 0 9568 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1667941163
transform 1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0692_
timestamp 1667941163
transform 1 0 13524 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0693_
timestamp 1667941163
transform 1 0 12972 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0694_
timestamp 1667941163
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0696_
timestamp 1667941163
transform 1 0 12604 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1667941163
transform 1 0 13800 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0698_
timestamp 1667941163
transform 1 0 14720 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0699_
timestamp 1667941163
transform 1 0 13156 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0700_
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0701_
timestamp 1667941163
transform 1 0 12052 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0702_
timestamp 1667941163
transform 1 0 11592 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0703_
timestamp 1667941163
transform 1 0 17664 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0705_
timestamp 1667941163
transform 1 0 13984 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 18952 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0707_
timestamp 1667941163
transform 1 0 17204 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0708_
timestamp 1667941163
transform 1 0 18216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _0709_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17756 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0710_
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_1  _0711_
timestamp 1667941163
transform 1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0712_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15824 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0713_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0714_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16192 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _0715_
timestamp 1667941163
transform 1 0 14812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0716_
timestamp 1667941163
transform 1 0 14996 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0717_
timestamp 1667941163
transform 1 0 14904 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _0718_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15088 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0719_
timestamp 1667941163
transform 1 0 15824 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0720_
timestamp 1667941163
transform 1 0 14444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0721_
timestamp 1667941163
transform 1 0 8372 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0722_
timestamp 1667941163
transform 1 0 7268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0723_
timestamp 1667941163
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0725_
timestamp 1667941163
transform 1 0 6164 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0726_
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0727_
timestamp 1667941163
transform 1 0 7452 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0728_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0729_
timestamp 1667941163
transform 1 0 7636 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0730_
timestamp 1667941163
transform 1 0 9108 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0731_
timestamp 1667941163
transform 1 0 8280 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0732_
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0733_
timestamp 1667941163
transform 1 0 8648 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0734_
timestamp 1667941163
transform 1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0735_
timestamp 1667941163
transform 1 0 9476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0736_
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0737_
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0738_
timestamp 1667941163
transform 1 0 5152 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0739_
timestamp 1667941163
transform 1 0 5060 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0740_
timestamp 1667941163
transform 1 0 7360 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0741_
timestamp 1667941163
transform 1 0 4876 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0742_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5520 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0743_
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0744_
timestamp 1667941163
transform 1 0 3312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0745_
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0746_
timestamp 1667941163
transform 1 0 5244 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0747_
timestamp 1667941163
transform 1 0 4140 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0748_
timestamp 1667941163
transform 1 0 3956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0749_
timestamp 1667941163
transform 1 0 4508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0750_
timestamp 1667941163
transform 1 0 4048 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0751_
timestamp 1667941163
transform 1 0 3864 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0752_
timestamp 1667941163
transform 1 0 3956 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0753_
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0754_
timestamp 1667941163
transform 1 0 4140 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0755_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4600 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0756_
timestamp 1667941163
transform 1 0 3956 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1667941163
transform 1 0 3220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0758_
timestamp 1667941163
transform 1 0 4416 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0760_
timestamp 1667941163
transform 1 0 4232 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0761_
timestamp 1667941163
transform 1 0 2576 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0762_
timestamp 1667941163
transform 1 0 5152 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0763_
timestamp 1667941163
transform 1 0 6072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0764_
timestamp 1667941163
transform 1 0 5520 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0765_
timestamp 1667941163
transform 1 0 5060 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0766_
timestamp 1667941163
transform 1 0 5796 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0767_
timestamp 1667941163
transform 1 0 6532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0768_
timestamp 1667941163
transform 1 0 6532 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 1667941163
transform 1 0 6532 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 5704 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0771_
timestamp 1667941163
transform 1 0 5796 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0772_
timestamp 1667941163
transform 1 0 5336 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0773_
timestamp 1667941163
transform 1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0774_
timestamp 1667941163
transform 1 0 6808 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0775_
timestamp 1667941163
transform 1 0 7636 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0776_
timestamp 1667941163
transform 1 0 7544 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1667941163
transform 1 0 7268 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1667941163
transform 1 0 8372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0779_
timestamp 1667941163
transform 1 0 9108 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1667941163
transform 1 0 8464 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0782_
timestamp 1667941163
transform 1 0 8004 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0783_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0784_
timestamp 1667941163
transform 1 0 9108 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0785_
timestamp 1667941163
transform 1 0 9016 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0786_
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0787_
timestamp 1667941163
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0788_
timestamp 1667941163
transform 1 0 6532 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0789_
timestamp 1667941163
transform 1 0 5336 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0790_
timestamp 1667941163
transform 1 0 5244 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0791_
timestamp 1667941163
transform 1 0 7728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0792_
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0793_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0794_
timestamp 1667941163
transform 1 0 6532 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0795_
timestamp 1667941163
transform 1 0 6440 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0796_
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0797_
timestamp 1667941163
transform 1 0 7912 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0798_
timestamp 1667941163
transform 1 0 5060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0799_
timestamp 1667941163
transform 1 0 4140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0800_
timestamp 1667941163
transform 1 0 3128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0801_
timestamp 1667941163
transform 1 0 5152 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0802_
timestamp 1667941163
transform 1 0 3128 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0803_
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0804_
timestamp 1667941163
transform 1 0 5612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0805_
timestamp 1667941163
transform 1 0 3128 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0806_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0807_
timestamp 1667941163
transform 1 0 2208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0809_
timestamp 1667941163
transform 1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0810_
timestamp 1667941163
transform 1 0 2392 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0811_
timestamp 1667941163
transform 1 0 2760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0812_
timestamp 1667941163
transform 1 0 3956 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0813_
timestamp 1667941163
transform 1 0 3404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0814_
timestamp 1667941163
transform 1 0 3220 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0815_
timestamp 1667941163
transform 1 0 4324 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0816_
timestamp 1667941163
transform 1 0 4232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0817_
timestamp 1667941163
transform 1 0 2944 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0819_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1667941163
transform 1 0 3220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0821_
timestamp 1667941163
transform 1 0 3864 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 3220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0823_
timestamp 1667941163
transform 1 0 3956 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1667941163
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0825_
timestamp 1667941163
transform 1 0 3956 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0826_
timestamp 1667941163
transform 1 0 3128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0827_
timestamp 1667941163
transform 1 0 4324 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0828_
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0829_
timestamp 1667941163
transform 1 0 4416 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0830_
timestamp 1667941163
transform 1 0 4968 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0831_
timestamp 1667941163
transform 1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0832_
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0833_
timestamp 1667941163
transform 1 0 5888 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0834_
timestamp 1667941163
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0835_
timestamp 1667941163
transform 1 0 4324 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0836_
timestamp 1667941163
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0837_
timestamp 1667941163
transform 1 0 6532 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0838_
timestamp 1667941163
transform 1 0 5520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0839_
timestamp 1667941163
transform 1 0 6256 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0840_
timestamp 1667941163
transform 1 0 8372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0841_
timestamp 1667941163
transform 1 0 6532 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0842_
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0843_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7268 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0844_
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0845_
timestamp 1667941163
transform 1 0 8096 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0846_
timestamp 1667941163
transform 1 0 7636 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0847_
timestamp 1667941163
transform 1 0 7636 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0848_
timestamp 1667941163
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0849_
timestamp 1667941163
transform 1 0 5888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0850_
timestamp 1667941163
transform 1 0 6532 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0851_
timestamp 1667941163
transform 1 0 6900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0852_
timestamp 1667941163
transform 1 0 5428 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0853_
timestamp 1667941163
transform 1 0 5520 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0854_
timestamp 1667941163
transform 1 0 6348 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0855_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6532 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0856_
timestamp 1667941163
transform 1 0 6532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 13616 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0859_
timestamp 1667941163
transform 1 0 13064 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0860_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0861_
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0862_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0863_
timestamp 1667941163
transform 1 0 12696 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0864_
timestamp 1667941163
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0865_
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0866_
timestamp 1667941163
transform 1 0 15272 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0867_
timestamp 1667941163
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0868_
timestamp 1667941163
transform 1 0 14812 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0870_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0871_
timestamp 1667941163
transform 1 0 13064 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0872_
timestamp 1667941163
transform 1 0 13248 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0873_
timestamp 1667941163
transform 1 0 13892 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0874_
timestamp 1667941163
transform 1 0 14904 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0875_
timestamp 1667941163
transform 1 0 8372 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0876_
timestamp 1667941163
transform 1 0 9108 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0877_
timestamp 1667941163
transform 1 0 9476 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0878_
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 1667941163
transform 1 0 10580 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0880_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0881_
timestamp 1667941163
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1667941163
transform 1 0 10396 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1667941163
transform 1 0 10212 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0884_
timestamp 1667941163
transform 1 0 10580 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0885_
timestamp 1667941163
transform 1 0 9292 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0886_
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0887_
timestamp 1667941163
transform 1 0 10948 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0888_
timestamp 1667941163
transform 1 0 10488 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0889_
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0890_
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0891_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0892_
timestamp 1667941163
transform 1 0 9568 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0893_
timestamp 1667941163
transform 1 0 9200 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1667941163
transform 1 0 12328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0895_
timestamp 1667941163
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0896_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0897_
timestamp 1667941163
transform 1 0 11960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0898_
timestamp 1667941163
transform 1 0 10672 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0899_
timestamp 1667941163
transform 1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0900_
timestamp 1667941163
transform 1 0 10672 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0901_
timestamp 1667941163
transform 1 0 8280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0902_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10396 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _0903_
timestamp 1667941163
transform 1 0 10212 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0904_
timestamp 1667941163
transform 1 0 9292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0905_
timestamp 1667941163
transform 1 0 8096 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1667941163
transform 1 0 13616 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1667941163
transform 1 0 11316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0909_
timestamp 1667941163
transform 1 0 13156 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0910_
timestamp 1667941163
transform 1 0 12144 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0911_
timestamp 1667941163
transform 1 0 13432 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0912_
timestamp 1667941163
transform 1 0 9384 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0913_
timestamp 1667941163
transform 1 0 9200 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1667941163
transform 1 0 10212 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 1667941163
transform 1 0 10304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0916_
timestamp 1667941163
transform 1 0 10304 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0917_
timestamp 1667941163
transform 1 0 12052 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0918_
timestamp 1667941163
transform 1 0 12696 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0919_
timestamp 1667941163
transform 1 0 11684 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0920_
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0921_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0922_
timestamp 1667941163
transform 1 0 11960 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0923_
timestamp 1667941163
transform 1 0 11684 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0924_
timestamp 1667941163
transform 1 0 9200 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0925_
timestamp 1667941163
transform 1 0 12236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0926_
timestamp 1667941163
transform 1 0 12512 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _0927_
timestamp 1667941163
transform 1 0 10120 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0928_
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0929_
timestamp 1667941163
transform 1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0930_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0931_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11316 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0932_
timestamp 1667941163
transform 1 0 9200 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1667941163
transform 1 0 10948 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0934_
timestamp 1667941163
transform 1 0 12328 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0935_
timestamp 1667941163
transform 1 0 12880 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _0936_
timestamp 1667941163
transform 1 0 9568 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0937_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0938_
timestamp 1667941163
transform 1 0 11684 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 1667941163
transform 1 0 12788 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0940_
timestamp 1667941163
transform 1 0 12696 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0941_
timestamp 1667941163
transform 1 0 22356 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0943_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0944_
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1667941163
transform 1 0 23000 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0946_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20976 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0947_
timestamp 1667941163
transform 1 0 21344 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0948_
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1667941163
transform 1 0 20056 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0950_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1667941163
transform 1 0 21896 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0952_
timestamp 1667941163
transform 1 0 20884 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0953_
timestamp 1667941163
transform 1 0 20516 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1667941163
transform 1 0 21712 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0955_
timestamp 1667941163
transform 1 0 19504 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1667941163
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0957_
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0958_
timestamp 1667941163
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0959_
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0960_
timestamp 1667941163
transform 1 0 20792 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0961_
timestamp 1667941163
transform 1 0 21068 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1667941163
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0963_
timestamp 1667941163
transform 1 0 20332 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0964_
timestamp 1667941163
transform 1 0 21160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0966_
timestamp 1667941163
transform 1 0 19412 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0967_
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0968_
timestamp 1667941163
transform 1 0 20148 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0969_
timestamp 1667941163
transform 1 0 17664 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0970_
timestamp 1667941163
transform 1 0 17664 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0972_
timestamp 1667941163
transform 1 0 16744 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0973_
timestamp 1667941163
transform 1 0 16376 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0974_
timestamp 1667941163
transform 1 0 14996 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0975_
timestamp 1667941163
transform 1 0 15364 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _0976_
timestamp 1667941163
transform 1 0 14904 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0977_
timestamp 1667941163
transform 1 0 13248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0978_
timestamp 1667941163
transform 1 0 15364 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0979_
timestamp 1667941163
transform 1 0 16376 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0980_
timestamp 1667941163
transform 1 0 17112 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0981_
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0982_
timestamp 1667941163
transform 1 0 16008 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0983_
timestamp 1667941163
transform 1 0 20700 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0984_
timestamp 1667941163
transform 1 0 18584 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0986_
timestamp 1667941163
transform 1 0 18952 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1667941163
transform 1 0 20424 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0988_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1667941163
transform 1 0 20056 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0990_
timestamp 1667941163
transform 1 0 19320 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0991_
timestamp 1667941163
transform 1 0 15272 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0992_
timestamp 1667941163
transform 1 0 16008 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0993_
timestamp 1667941163
transform 1 0 15732 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 16100 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0995_
timestamp 1667941163
transform 1 0 16836 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0996_
timestamp 1667941163
transform 1 0 15824 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1667941163
transform 1 0 15916 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0998_
timestamp 1667941163
transform 1 0 14352 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0999_
timestamp 1667941163
transform 1 0 13432 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1000_
timestamp 1667941163
transform 1 0 15456 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1001_
timestamp 1667941163
transform 1 0 14536 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1002_
timestamp 1667941163
transform 1 0 16100 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 17664 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1004_
timestamp 1667941163
transform 1 0 15272 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1005_
timestamp 1667941163
transform 1 0 14260 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1006_
timestamp 1667941163
transform 1 0 14444 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 14260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1008_
timestamp 1667941163
transform 1 0 14260 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1009_
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1010_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1011_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10580 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1667941163
transform 1 0 17940 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1667941163
transform 1 0 19780 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1667941163
transform 1 0 20056 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1667941163
transform 1 0 22080 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1667941163
transform 1 0 18492 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1667941163
transform 1 0 12420 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1667941163
transform 1 0 8372 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1667941163
transform 1 0 9476 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1667941163
transform 1 0 17112 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1667941163
transform 1 0 15640 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1667941163
transform 1 0 6532 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1667941163
transform 1 0 9476 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1667941163
transform 1 0 2116 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1667941163
transform 1 0 2392 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1667941163
transform 1 0 6532 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1667941163
transform 1 0 9568 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1667941163
transform 1 0 4600 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1667941163
transform 1 0 8004 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1667941163
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1667941163
transform 1 0 8740 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1667941163
transform 1 0 6992 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1667941163
transform 1 0 6532 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1667941163
transform 1 0 8372 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1667941163
transform 1 0 9752 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1667941163
transform 1 0 11316 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1046_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12144 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1667941163
transform 1 0 22448 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1667941163
transform 1 0 22172 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1667941163
transform 1 0 22080 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1667941163
transform 1 0 21988 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1667941163
transform 1 0 21160 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1667941163
transform 1 0 19320 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1667941163
transform 1 0 16928 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1667941163
transform 1 0 17480 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1062_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1667941163
transform 1 0 16008 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1667941163
transform 1 0 13984 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1667941163
transform 1 0 16652 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1667941163
transform 1 0 14904 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1667941163
transform 1 0 13248 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1071_
timestamp 1667941163
transform 1 0 37352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1667941163
transform 1 0 37812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1073_
timestamp 1667941163
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1667941163
transform 1 0 2300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1667941163
transform 1 0 9016 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout24 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout26
timestamp 1667941163
transform 1 0 6348 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout27
timestamp 1667941163
transform 1 0 2392 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout28
timestamp 1667941163
transform 1 0 10304 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout29
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout30
timestamp 1667941163
transform 1 0 2576 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout31
timestamp 1667941163
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout32
timestamp 1667941163
transform 1 0 17572 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout33
timestamp 1667941163
transform 1 0 18676 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout34
timestamp 1667941163
transform 1 0 13524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout36
timestamp 1667941163
transform 1 0 13524 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1667941163
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout38
timestamp 1667941163
transform 1 0 12328 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout39
timestamp 1667941163
transform 1 0 3772 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1667941163
transform 1 0 37444 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 38088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1667941163
transform 1 0 32936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1667941163
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  solo_squash_caravel_40 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38088 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  solo_squash_caravel_41
timestamp 1667941163
transform 1 0 38088 0 -1 19584
box -38 -48 314 592
<< labels >>
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 blue
port 0 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 debug_design_reset
port 1 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 debug_gpio_ready
port 2 nsew signal tristate
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 debug_oeb[0]
port 3 nsew signal tristate
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 debug_oeb[1]
port 4 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 design_oeb[0]
port 5 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 design_oeb[1]
port 6 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 design_oeb[2]
port 7 nsew signal tristate
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 design_oeb[3]
port 8 nsew signal tristate
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 design_oeb[4]
port 9 nsew signal tristate
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 design_oeb[5]
port 10 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 down_key_n
port 11 nsew signal input
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 ext_reset_n
port 12 nsew signal input
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 gpio_ready
port 13 nsew signal input
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 green
port 14 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 hsync
port 15 nsew signal tristate
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 new_game_n
port 16 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 pause_n
port 17 nsew signal input
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 red
port 18 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 speaker
port 19 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 up_key_n
port 20 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 22 nsew ground bidirectional
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 vsync
port 23 nsew signal tristate
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 wb_clk_i
port 24 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 wb_rst_i
port 25 nsew signal input
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 10800 28526 10800 28526 0 _0000_
rlabel metal2 17894 31110 17894 31110 0 _0001_
rlabel metal1 19964 31654 19964 31654 0 _0002_
rlabel via1 20373 30226 20373 30226 0 _0003_
rlabel metal1 22346 26350 22346 26350 0 _0004_
rlabel metal2 18354 16966 18354 16966 0 _0005_
rlabel metal1 9701 16558 9701 16558 0 _0006_
rlabel viali 12727 17170 12727 17170 0 _0007_
rlabel metal2 9154 14790 9154 14790 0 _0008_
rlabel metal2 9982 13090 9982 13090 0 _0009_
rlabel metal1 12128 13226 12128 13226 0 _0010_
rlabel metal2 17986 14994 17986 14994 0 _0011_
rlabel metal1 17332 13906 17332 13906 0 _0012_
rlabel via1 15957 13294 15957 13294 0 _0013_
rlabel metal2 6210 26758 6210 26758 0 _0014_
rlabel metal1 9660 25738 9660 25738 0 _0015_
rlabel metal1 2433 26282 2433 26282 0 _0016_
rlabel metal1 2484 27642 2484 27642 0 _0017_
rlabel metal1 2668 29818 2668 29818 0 _0018_
rlabel via1 6849 32402 6849 32402 0 _0019_
rlabel metal1 8372 32538 8372 32538 0 _0020_
rlabel metal1 9782 33558 9782 33558 0 _0021_
rlabel metal1 5101 24854 5101 24854 0 _0022_
rlabel metal1 8132 24786 8132 24786 0 _0023_
rlabel metal1 2065 24174 2065 24174 0 _0024_
rlabel metal1 4768 21930 4768 21930 0 _0025_
rlabel metal1 2019 19822 2019 19822 0 _0026_
rlabel metal2 4094 16966 4094 16966 0 _0027_
rlabel metal1 8724 18326 8724 18326 0 _0028_
rlabel metal1 7268 16218 7268 16218 0 _0029_
rlabel metal1 6700 22678 6700 22678 0 _0030_
rlabel metal2 14950 23970 14950 23970 0 _0031_
rlabel metal1 8648 23290 8648 23290 0 _0032_
rlabel metal1 10713 27030 10713 27030 0 _0033_
rlabel metal2 12190 23970 12190 23970 0 _0034_
rlabel metal2 12742 32674 12742 32674 0 _0035_
rlabel metal2 23046 21318 23046 21318 0 _0036_
rlabel metal1 21528 22202 21528 22202 0 _0037_
rlabel metal1 22011 22950 22011 22950 0 _0038_
rlabel metal2 22126 24514 22126 24514 0 _0039_
rlabel metal1 19258 21930 19258 21930 0 _0040_
rlabel metal1 17567 21522 17567 21522 0 _0041_
rlabel metal1 22535 19822 22535 19822 0 _0042_
rlabel metal1 21753 18734 21753 18734 0 _0043_
rlabel metal1 19959 18326 19959 18326 0 _0044_
rlabel metal2 17710 19346 17710 19346 0 _0045_
rlabel metal1 14352 22066 14352 22066 0 _0046_
rlabel metal2 17158 22882 17158 22882 0 _0047_
rlabel metal1 16330 23562 16330 23562 0 _0048_
rlabel metal2 18998 26486 18998 26486 0 _0049_
rlabel metal2 19366 25007 19366 25007 0 _0050_
rlabel metal1 17056 30226 17056 30226 0 _0051_
rlabel metal1 16228 32878 16228 32878 0 _0052_
rlabel metal1 13662 32266 13662 32266 0 _0053_
rlabel metal1 17337 31790 17337 31790 0 _0054_
rlabel metal1 14750 29206 14750 29206 0 _0055_
rlabel metal1 14163 28118 14163 28118 0 _0056_
rlabel metal1 17572 18258 17572 18258 0 _0057_
rlabel metal1 17434 19346 17434 19346 0 _0058_
rlabel via1 16330 18870 16330 18870 0 _0059_
rlabel via1 18170 18717 18170 18717 0 _0060_
rlabel metal1 19918 19788 19918 19788 0 _0061_
rlabel metal1 15962 20026 15962 20026 0 _0062_
rlabel metal1 15870 19822 15870 19822 0 _0063_
rlabel metal2 17526 25772 17526 25772 0 _0064_
rlabel metal1 18216 26894 18216 26894 0 _0065_
rlabel metal2 12926 26078 12926 26078 0 _0066_
rlabel metal1 17618 25670 17618 25670 0 _0067_
rlabel metal1 13984 19754 13984 19754 0 _0068_
rlabel metal1 17526 25262 17526 25262 0 _0069_
rlabel metal2 17894 25092 17894 25092 0 _0070_
rlabel metal1 18538 24752 18538 24752 0 _0071_
rlabel metal1 19412 23154 19412 23154 0 _0072_
rlabel metal1 17664 24310 17664 24310 0 _0073_
rlabel metal1 20884 21590 20884 21590 0 _0074_
rlabel metal1 19734 23290 19734 23290 0 _0075_
rlabel metal2 21850 21760 21850 21760 0 _0076_
rlabel metal1 20056 24174 20056 24174 0 _0077_
rlabel metal2 19734 24514 19734 24514 0 _0078_
rlabel via2 14858 27421 14858 27421 0 _0079_
rlabel metal1 11362 31790 11362 31790 0 _0080_
rlabel metal2 13662 27234 13662 27234 0 _0081_
rlabel metal2 14858 22678 14858 22678 0 _0082_
rlabel metal1 13754 20570 13754 20570 0 _0083_
rlabel metal1 14858 26826 14858 26826 0 _0084_
rlabel metal1 13202 26758 13202 26758 0 _0085_
rlabel metal1 14628 24718 14628 24718 0 _0086_
rlabel metal1 15732 24786 15732 24786 0 _0087_
rlabel metal1 9430 32436 9430 32436 0 _0088_
rlabel metal1 9522 31960 9522 31960 0 _0089_
rlabel metal1 13915 32198 13915 32198 0 _0090_
rlabel metal2 14490 29750 14490 29750 0 _0091_
rlabel metal1 23230 24616 23230 24616 0 _0092_
rlabel metal1 15502 24922 15502 24922 0 _0093_
rlabel metal2 20746 25024 20746 25024 0 _0094_
rlabel metal1 14674 26350 14674 26350 0 _0095_
rlabel metal2 17158 27166 17158 27166 0 _0096_
rlabel metal1 14490 26248 14490 26248 0 _0097_
rlabel via2 2070 26979 2070 26979 0 _0098_
rlabel metal1 12972 21114 12972 21114 0 _0099_
rlabel metal2 20378 20128 20378 20128 0 _0100_
rlabel metal1 19182 19890 19182 19890 0 _0101_
rlabel metal2 19458 20026 19458 20026 0 _0102_
rlabel metal1 19872 14382 19872 14382 0 _0103_
rlabel metal1 13570 19380 13570 19380 0 _0104_
rlabel metal1 24748 26962 24748 26962 0 _0105_
rlabel metal1 24380 27098 24380 27098 0 _0106_
rlabel metal1 22172 29138 22172 29138 0 _0107_
rlabel metal1 18860 28390 18860 28390 0 _0108_
rlabel metal2 18814 28254 18814 28254 0 _0109_
rlabel metal2 18998 28356 18998 28356 0 _0110_
rlabel metal1 19412 28594 19412 28594 0 _0111_
rlabel metal1 21114 28594 21114 28594 0 _0112_
rlabel metal1 20470 28084 20470 28084 0 _0113_
rlabel metal1 24334 28016 24334 28016 0 _0114_
rlabel metal1 24472 28118 24472 28118 0 _0115_
rlabel metal1 24426 27438 24426 27438 0 _0116_
rlabel metal1 23966 26010 23966 26010 0 _0117_
rlabel metal2 22402 28730 22402 28730 0 _0118_
rlabel metal1 22908 31450 22908 31450 0 _0119_
rlabel metal1 23184 29818 23184 29818 0 _0120_
rlabel metal1 22816 30362 22816 30362 0 _0121_
rlabel metal1 23184 28526 23184 28526 0 _0122_
rlabel metal1 22310 28186 22310 28186 0 _0123_
rlabel metal1 23092 29138 23092 29138 0 _0124_
rlabel metal2 24978 26520 24978 26520 0 _0125_
rlabel metal2 24794 26554 24794 26554 0 _0126_
rlabel metal1 18078 27370 18078 27370 0 _0127_
rlabel metal1 24702 26486 24702 26486 0 _0128_
rlabel metal2 25070 27030 25070 27030 0 _0129_
rlabel metal1 24978 29546 24978 29546 0 _0130_
rlabel metal1 23000 30226 23000 30226 0 _0131_
rlabel metal1 24242 30838 24242 30838 0 _0132_
rlabel metal1 24748 30702 24748 30702 0 _0133_
rlabel metal1 24656 30906 24656 30906 0 _0134_
rlabel metal2 20746 28084 20746 28084 0 _0135_
rlabel metal2 22954 28866 22954 28866 0 _0136_
rlabel metal1 23414 29070 23414 29070 0 _0137_
rlabel metal1 23092 25466 23092 25466 0 _0138_
rlabel metal1 24702 28628 24702 28628 0 _0139_
rlabel metal2 25070 28900 25070 28900 0 _0140_
rlabel metal2 25070 29444 25070 29444 0 _0141_
rlabel metal1 24610 31280 24610 31280 0 _0142_
rlabel metal2 25346 30838 25346 30838 0 _0143_
rlabel metal1 9522 31790 9522 31790 0 _0144_
rlabel metal1 6302 31450 6302 31450 0 _0145_
rlabel metal1 8924 31994 8924 31994 0 _0146_
rlabel metal2 11086 32640 11086 32640 0 _0147_
rlabel metal2 7774 30906 7774 30906 0 _0148_
rlabel metal2 4186 28237 4186 28237 0 _0149_
rlabel metal1 9706 30736 9706 30736 0 _0150_
rlabel metal2 8050 30906 8050 30906 0 _0151_
rlabel metal1 8418 18904 8418 18904 0 _0152_
rlabel metal1 8510 22032 8510 22032 0 _0153_
rlabel metal2 12374 21488 12374 21488 0 _0154_
rlabel metal1 5382 18326 5382 18326 0 _0155_
rlabel metal2 7958 21250 7958 21250 0 _0156_
rlabel metal1 7774 30634 7774 30634 0 _0157_
rlabel metal2 14490 31416 14490 31416 0 _0158_
rlabel metal1 14582 32878 14582 32878 0 _0159_
rlabel metal2 20562 23936 20562 23936 0 _0160_
rlabel metal1 15640 20434 15640 20434 0 _0161_
rlabel metal1 15088 20230 15088 20230 0 _0162_
rlabel metal2 18354 27608 18354 27608 0 _0163_
rlabel metal1 15686 27574 15686 27574 0 _0164_
rlabel metal1 14996 26962 14996 26962 0 _0165_
rlabel metal2 14398 25262 14398 25262 0 _0166_
rlabel via2 14950 25109 14950 25109 0 _0167_
rlabel metal2 5888 18666 5888 18666 0 _0168_
rlabel metal1 16238 19482 16238 19482 0 _0169_
rlabel metal1 17204 27030 17204 27030 0 _0170_
rlabel metal1 16200 26282 16200 26282 0 _0171_
rlabel metal1 16652 26350 16652 26350 0 _0172_
rlabel metal1 16468 17170 16468 17170 0 _0173_
rlabel metal1 11316 29274 11316 29274 0 _0174_
rlabel metal1 18446 18326 18446 18326 0 _0175_
rlabel metal1 13064 21998 13064 21998 0 _0176_
rlabel metal2 20562 29308 20562 29308 0 _0177_
rlabel metal1 16422 17034 16422 17034 0 _0178_
rlabel metal2 17894 29376 17894 29376 0 _0179_
rlabel metal2 18446 30260 18446 30260 0 _0180_
rlabel metal1 19274 30906 19274 30906 0 _0181_
rlabel metal1 18860 30362 18860 30362 0 _0182_
rlabel metal1 19458 30838 19458 30838 0 _0183_
rlabel metal1 21482 29478 21482 29478 0 _0184_
rlabel metal2 20102 29376 20102 29376 0 _0185_
rlabel metal1 20516 29818 20516 29818 0 _0186_
rlabel metal2 22126 27132 22126 27132 0 _0187_
rlabel metal1 12926 18326 12926 18326 0 _0188_
rlabel metal1 16882 27370 16882 27370 0 _0189_
rlabel metal2 15410 26826 15410 26826 0 _0190_
rlabel via2 15594 16643 15594 16643 0 _0191_
rlabel metal2 15594 13362 15594 13362 0 _0192_
rlabel metal1 16008 15606 16008 15606 0 _0193_
rlabel metal2 18630 13634 18630 13634 0 _0194_
rlabel metal1 16560 14246 16560 14246 0 _0195_
rlabel metal2 15778 15844 15778 15844 0 _0196_
rlabel metal2 16146 17204 16146 17204 0 _0197_
rlabel metal1 12788 18054 12788 18054 0 _0198_
rlabel metal1 18676 16558 18676 16558 0 _0199_
rlabel metal1 8234 32980 8234 32980 0 _0200_
rlabel metal1 10442 17646 10442 17646 0 _0201_
rlabel metal2 9890 13974 9890 13974 0 _0202_
rlabel metal1 13685 19822 13685 19822 0 _0203_
rlabel metal1 9338 17204 9338 17204 0 _0204_
rlabel metal1 9844 17170 9844 17170 0 _0205_
rlabel metal1 10672 16082 10672 16082 0 _0206_
rlabel metal2 14766 25551 14766 25551 0 _0207_
rlabel metal1 6854 21080 6854 21080 0 _0208_
rlabel metal1 15088 14042 15088 14042 0 _0209_
rlabel metal2 11822 16014 11822 16014 0 _0210_
rlabel metal2 13754 13532 13754 13532 0 _0211_
rlabel metal1 11822 16660 11822 16660 0 _0212_
rlabel metal2 11178 17000 11178 17000 0 _0213_
rlabel metal1 11546 17102 11546 17102 0 _0214_
rlabel metal2 11730 17782 11730 17782 0 _0215_
rlabel metal1 12742 17850 12742 17850 0 _0216_
rlabel metal2 12742 16320 12742 16320 0 _0217_
rlabel metal1 11546 14348 11546 14348 0 _0218_
rlabel metal2 13018 15436 13018 15436 0 _0219_
rlabel metal1 12052 14586 12052 14586 0 _0220_
rlabel metal1 11638 15674 11638 15674 0 _0221_
rlabel metal1 10166 15980 10166 15980 0 _0222_
rlabel metal1 11316 14994 11316 14994 0 _0223_
rlabel metal2 12650 14314 12650 14314 0 _0224_
rlabel metal1 9154 14416 9154 14416 0 _0225_
rlabel metal1 11500 13838 11500 13838 0 _0226_
rlabel metal2 10810 13260 10810 13260 0 _0227_
rlabel metal2 10902 13464 10902 13464 0 _0228_
rlabel metal2 9890 13260 9890 13260 0 _0229_
rlabel metal1 13294 17680 13294 17680 0 _0230_
rlabel metal1 13800 14994 13800 14994 0 _0231_
rlabel metal1 12788 14586 12788 14586 0 _0232_
rlabel metal1 13800 14586 13800 14586 0 _0233_
rlabel metal1 13248 12818 13248 12818 0 _0234_
rlabel metal2 14766 13090 14766 13090 0 _0235_
rlabel metal2 14398 13940 14398 13940 0 _0236_
rlabel metal1 13386 12954 13386 12954 0 _0237_
rlabel metal1 12972 13906 12972 13906 0 _0238_
rlabel metal2 11638 13498 11638 13498 0 _0239_
rlabel metal1 17894 14926 17894 14926 0 _0240_
rlabel metal2 14490 14790 14490 14790 0 _0241_
rlabel metal1 15962 14518 15962 14518 0 _0242_
rlabel metal1 17618 16660 17618 16660 0 _0243_
rlabel metal2 18078 15538 18078 15538 0 _0244_
rlabel metal1 19458 18394 19458 18394 0 _0245_
rlabel metal1 18814 16014 18814 16014 0 _0246_
rlabel metal1 15548 15674 15548 15674 0 _0247_
rlabel metal1 17204 15538 17204 15538 0 _0248_
rlabel metal1 17388 15334 17388 15334 0 _0249_
rlabel metal2 15318 16422 15318 16422 0 _0250_
rlabel metal1 15088 15130 15088 15130 0 _0251_
rlabel metal2 15318 17051 15318 17051 0 _0252_
rlabel metal1 14674 17136 14674 17136 0 _0253_
rlabel metal2 14490 17476 14490 17476 0 _0254_
rlabel metal2 12098 26078 12098 26078 0 _0255_
rlabel metal1 6486 19754 6486 19754 0 _0256_
rlabel metal1 4692 20026 4692 20026 0 _0257_
rlabel metal1 6670 26384 6670 26384 0 _0258_
rlabel metal2 7590 25466 7590 25466 0 _0259_
rlabel metal1 4186 26248 4186 26248 0 _0260_
rlabel metal1 9476 25466 9476 25466 0 _0261_
rlabel metal1 7912 26282 7912 26282 0 _0262_
rlabel metal1 9062 27438 9062 27438 0 _0263_
rlabel metal2 8326 26622 8326 26622 0 _0264_
rlabel metal2 8602 25670 8602 25670 0 _0265_
rlabel metal1 9798 25840 9798 25840 0 _0266_
rlabel metal1 12788 23698 12788 23698 0 _0267_
rlabel metal2 2346 21318 2346 21318 0 _0268_
rlabel metal1 5796 28526 5796 28526 0 _0269_
rlabel metal2 5290 26452 5290 26452 0 _0270_
rlabel metal1 5750 25840 5750 25840 0 _0271_
rlabel metal2 5566 26180 5566 26180 0 _0272_
rlabel metal2 4922 26214 4922 26214 0 _0273_
rlabel metal1 4884 26010 4884 26010 0 _0274_
rlabel metal1 5060 25738 5060 25738 0 _0275_
rlabel metal1 2530 25908 2530 25908 0 _0276_
rlabel metal1 4738 28050 4738 28050 0 _0277_
rlabel metal2 4002 28220 4002 28220 0 _0278_
rlabel metal1 4524 27030 4524 27030 0 _0279_
rlabel metal2 4094 25670 4094 25670 0 _0280_
rlabel metal1 4232 25942 4232 25942 0 _0281_
rlabel metal1 4462 26010 4462 26010 0 _0282_
rlabel metal1 2530 27404 2530 27404 0 _0283_
rlabel metal1 4508 27642 4508 27642 0 _0284_
rlabel metal1 5612 29682 5612 29682 0 _0285_
rlabel metal1 3910 29478 3910 29478 0 _0286_
rlabel metal1 4248 30226 4248 30226 0 _0287_
rlabel metal2 4462 30464 4462 30464 0 _0288_
rlabel metal1 9890 32402 9890 32402 0 _0289_
rlabel metal1 2622 29648 2622 29648 0 _0290_
rlabel metal1 5796 31926 5796 31926 0 _0291_
rlabel metal2 9430 27846 9430 27846 0 _0292_
rlabel metal1 5842 30634 5842 30634 0 _0293_
rlabel metal1 5842 30770 5842 30770 0 _0294_
rlabel metal1 6348 30634 6348 30634 0 _0295_
rlabel metal2 6670 30532 6670 30532 0 _0296_
rlabel metal1 7084 29274 7084 29274 0 _0297_
rlabel metal1 5704 28186 5704 28186 0 _0298_
rlabel metal1 5888 29682 5888 29682 0 _0299_
rlabel metal1 6900 28526 6900 28526 0 _0300_
rlabel metal1 8556 29138 8556 29138 0 _0301_
rlabel metal1 7498 28594 7498 28594 0 _0302_
rlabel metal2 8050 28356 8050 28356 0 _0303_
rlabel metal1 7544 28730 7544 28730 0 _0304_
rlabel metal1 8142 32402 8142 32402 0 _0305_
rlabel metal1 9568 29614 9568 29614 0 _0306_
rlabel metal1 8924 29478 8924 29478 0 _0307_
rlabel metal1 8050 29104 8050 29104 0 _0308_
rlabel metal1 9338 29036 9338 29036 0 _0309_
rlabel metal1 9384 29138 9384 29138 0 _0310_
rlabel metal2 9522 28628 9522 28628 0 _0311_
rlabel metal1 8740 29274 8740 29274 0 _0312_
rlabel metal1 9246 33082 9246 33082 0 _0313_
rlabel metal2 9982 25024 9982 25024 0 _0314_
rlabel metal1 5750 22746 5750 22746 0 _0315_
rlabel metal1 8050 23834 8050 23834 0 _0316_
rlabel metal1 6716 25466 6716 25466 0 _0317_
rlabel metal2 6118 24004 6118 24004 0 _0318_
rlabel metal1 7084 24378 7084 24378 0 _0319_
rlabel metal2 7130 24650 7130 24650 0 _0320_
rlabel metal1 7866 24174 7866 24174 0 _0321_
rlabel metal1 2530 21998 2530 21998 0 _0322_
rlabel metal1 3404 21930 3404 21930 0 _0323_
rlabel metal1 5566 20468 5566 20468 0 _0324_
rlabel metal1 2622 21488 2622 21488 0 _0325_
rlabel metal1 2530 23732 2530 23732 0 _0326_
rlabel metal1 3358 23664 3358 23664 0 _0327_
rlabel metal2 3450 23970 3450 23970 0 _0328_
rlabel metal1 4186 23630 4186 23630 0 _0329_
rlabel metal2 2346 24582 2346 24582 0 _0330_
rlabel metal2 2162 21794 2162 21794 0 _0331_
rlabel metal1 2990 21964 2990 21964 0 _0332_
rlabel metal2 2806 22134 2806 22134 0 _0333_
rlabel metal1 3174 21522 3174 21522 0 _0334_
rlabel metal2 3450 22814 3450 22814 0 _0335_
rlabel metal1 3404 22406 3404 22406 0 _0336_
rlabel metal1 4186 21522 4186 21522 0 _0337_
rlabel metal1 4324 21658 4324 21658 0 _0338_
rlabel metal1 4186 20366 4186 20366 0 _0339_
rlabel metal1 3726 22066 3726 22066 0 _0340_
rlabel metal2 3266 21386 3266 21386 0 _0341_
rlabel metal2 3450 20570 3450 20570 0 _0342_
rlabel metal1 4140 19686 4140 19686 0 _0343_
rlabel metal2 12006 20060 12006 20060 0 _0344_
rlabel metal2 2254 20230 2254 20230 0 _0345_
rlabel metal2 4462 18445 4462 18445 0 _0346_
rlabel metal2 3082 19244 3082 19244 0 _0347_
rlabel metal2 4646 18428 4646 18428 0 _0348_
rlabel metal1 4002 18326 4002 18326 0 _0349_
rlabel metal1 4922 17646 4922 17646 0 _0350_
rlabel metal1 4830 16558 4830 16558 0 _0351_
rlabel metal1 8740 18938 8740 18938 0 _0352_
rlabel metal1 6624 18326 6624 18326 0 _0353_
rlabel metal1 4324 18394 4324 18394 0 _0354_
rlabel metal2 5566 18972 5566 18972 0 _0355_
rlabel metal1 6118 19346 6118 19346 0 _0356_
rlabel metal1 6716 18938 6716 18938 0 _0357_
rlabel metal1 6172 18598 6172 18598 0 _0358_
rlabel metal1 6670 18632 6670 18632 0 _0359_
rlabel metal2 7130 17952 7130 17952 0 _0360_
rlabel metal1 7728 18802 7728 18802 0 _0361_
rlabel metal1 7866 17850 7866 17850 0 _0362_
rlabel metal2 7866 18428 7866 18428 0 _0363_
rlabel metal1 8326 18258 8326 18258 0 _0364_
rlabel metal2 7866 17612 7866 17612 0 _0365_
rlabel metal2 7406 16524 7406 16524 0 _0366_
rlabel metal1 6440 22950 6440 22950 0 _0367_
rlabel metal1 6348 20026 6348 20026 0 _0368_
rlabel metal1 6440 20570 6440 20570 0 _0369_
rlabel metal1 6210 20910 6210 20910 0 _0370_
rlabel metal1 6210 20978 6210 20978 0 _0371_
rlabel metal1 6716 20026 6716 20026 0 _0372_
rlabel metal1 6992 23086 6992 23086 0 _0373_
rlabel metal2 13478 17952 13478 17952 0 _0374_
rlabel via1 13570 18258 13570 18258 0 _0375_
rlabel metal1 13202 17850 13202 17850 0 _0376_
rlabel metal1 13984 18938 13984 18938 0 _0377_
rlabel metal2 17986 17986 17986 17986 0 _0378_
rlabel metal2 14122 18564 14122 18564 0 _0379_
rlabel metal2 13110 20026 13110 20026 0 _0380_
rlabel metal2 14306 19176 14306 19176 0 _0381_
rlabel metal1 15594 21522 15594 21522 0 _0382_
rlabel metal1 16882 21930 16882 21930 0 _0383_
rlabel metal1 16560 21658 16560 21658 0 _0384_
rlabel metal1 15318 18224 15318 18224 0 _0385_
rlabel metal1 16284 21114 16284 21114 0 _0386_
rlabel metal1 14858 21930 14858 21930 0 _0387_
rlabel metal2 13478 24650 13478 24650 0 _0388_
rlabel metal1 13800 23494 13800 23494 0 _0389_
rlabel metal1 14812 23698 14812 23698 0 _0390_
rlabel metal1 8280 23018 8280 23018 0 _0391_
rlabel metal1 9522 21114 9522 21114 0 _0392_
rlabel metal2 10994 20128 10994 20128 0 _0393_
rlabel metal1 9200 21998 9200 21998 0 _0394_
rlabel metal1 10764 24854 10764 24854 0 _0395_
rlabel metal1 10626 24752 10626 24752 0 _0396_
rlabel metal1 10304 24854 10304 24854 0 _0397_
rlabel metal1 10534 24378 10534 24378 0 _0398_
rlabel metal1 11408 21522 11408 21522 0 _0399_
rlabel via1 11178 22678 11178 22678 0 _0400_
rlabel metal1 11132 21930 11132 21930 0 _0401_
rlabel metal1 10994 21352 10994 21352 0 _0402_
rlabel metal2 11914 21454 11914 21454 0 _0403_
rlabel metal1 11224 20910 11224 20910 0 _0404_
rlabel metal1 12006 22202 12006 22202 0 _0405_
rlabel metal2 12742 22372 12742 22372 0 _0406_
rlabel metal1 10580 22066 10580 22066 0 _0407_
rlabel metal2 9614 22644 9614 22644 0 _0408_
rlabel metal1 10120 22610 10120 22610 0 _0409_
rlabel metal2 11730 20672 11730 20672 0 _0410_
rlabel metal2 12190 20604 12190 20604 0 _0411_
rlabel metal1 11638 20570 11638 20570 0 _0412_
rlabel metal1 11546 20026 11546 20026 0 _0413_
rlabel metal1 10764 20570 10764 20570 0 _0414_
rlabel metal2 10902 20366 10902 20366 0 _0415_
rlabel metal1 10994 21114 10994 21114 0 _0416_
rlabel metal1 9522 21046 9522 21046 0 _0417_
rlabel metal1 10534 21114 10534 21114 0 _0418_
rlabel metal2 10258 22882 10258 22882 0 _0419_
rlabel metal1 8878 23222 8878 23222 0 _0420_
rlabel metal2 12098 27200 12098 27200 0 _0421_
rlabel metal2 12006 27268 12006 27268 0 _0422_
rlabel metal1 12374 23732 12374 23732 0 _0423_
rlabel metal2 16422 23630 16422 23630 0 _0424_
rlabel metal1 10120 31858 10120 31858 0 _0425_
rlabel metal2 9936 31314 9936 31314 0 _0426_
rlabel metal2 10626 31994 10626 31994 0 _0427_
rlabel metal2 10718 31008 10718 31008 0 _0428_
rlabel metal1 10994 31790 10994 31790 0 _0429_
rlabel metal2 12466 26656 12466 26656 0 _0430_
rlabel metal2 13110 26996 13110 26996 0 _0431_
rlabel metal2 12282 26962 12282 26962 0 _0432_
rlabel metal1 12328 27574 12328 27574 0 _0433_
rlabel metal2 12282 29580 12282 29580 0 _0434_
rlabel metal2 12558 29954 12558 29954 0 _0435_
rlabel metal1 12098 32198 12098 32198 0 _0436_
rlabel metal1 9292 30702 9292 30702 0 _0437_
rlabel metal1 13064 30362 13064 30362 0 _0438_
rlabel metal1 12788 30906 12788 30906 0 _0439_
rlabel metal2 10626 31042 10626 31042 0 _0440_
rlabel metal1 10902 32368 10902 32368 0 _0441_
rlabel metal1 11638 31824 11638 31824 0 _0442_
rlabel metal1 12282 31382 12282 31382 0 _0443_
rlabel metal2 11362 31382 11362 31382 0 _0444_
rlabel metal2 9890 30719 9890 30719 0 _0445_
rlabel metal2 12650 29614 12650 29614 0 _0446_
rlabel metal2 13294 30328 13294 30328 0 _0447_
rlabel metal1 12650 31246 12650 31246 0 _0448_
rlabel metal1 11178 30770 11178 30770 0 _0449_
rlabel metal2 11914 31110 11914 31110 0 _0450_
rlabel metal2 12466 31552 12466 31552 0 _0451_
rlabel metal2 13202 32198 13202 32198 0 _0452_
rlabel metal2 21758 21794 21758 21794 0 _0453_
rlabel metal1 17710 19244 17710 19244 0 _0454_
rlabel metal2 18998 19210 18998 19210 0 _0455_
rlabel metal1 22908 20910 22908 20910 0 _0456_
rlabel metal1 21390 22406 21390 22406 0 _0457_
rlabel metal1 21574 21658 21574 21658 0 _0458_
rlabel metal1 20424 22746 20424 22746 0 _0459_
rlabel metal1 22264 23086 22264 23086 0 _0460_
rlabel metal2 20930 23834 20930 23834 0 _0461_
rlabel metal1 21528 24174 21528 24174 0 _0462_
rlabel metal1 19228 21114 19228 21114 0 _0463_
rlabel metal1 18262 20842 18262 20842 0 _0464_
rlabel metal1 21206 20026 21206 20026 0 _0465_
rlabel metal1 21160 20570 21160 20570 0 _0466_
rlabel metal2 22954 20604 22954 20604 0 _0467_
rlabel metal1 19228 19210 19228 19210 0 _0468_
rlabel metal1 21758 19346 21758 19346 0 _0469_
rlabel metal1 20102 19142 20102 19142 0 _0470_
rlabel metal2 20194 19074 20194 19074 0 _0471_
rlabel metal1 17940 18734 17940 18734 0 _0472_
rlabel metal1 17434 16218 17434 16218 0 _0473_
rlabel metal1 17204 21862 17204 21862 0 _0474_
rlabel metal2 15226 17476 15226 17476 0 _0475_
rlabel metal1 15502 18190 15502 18190 0 _0476_
rlabel metal1 15364 21114 15364 21114 0 _0477_
rlabel metal1 14306 21658 14306 21658 0 _0478_
rlabel metal1 19464 24752 19464 24752 0 _0479_
rlabel metal2 16330 23647 16330 23647 0 _0480_
rlabel metal1 16192 23290 16192 23290 0 _0481_
rlabel metal1 19780 26350 19780 26350 0 _0482_
rlabel metal1 18630 25364 18630 25364 0 _0483_
rlabel metal2 19182 25670 19182 25670 0 _0484_
rlabel metal1 20424 24922 20424 24922 0 _0485_
rlabel metal1 19964 26418 19964 26418 0 _0486_
rlabel metal1 19550 24854 19550 24854 0 _0487_
rlabel metal1 15870 33286 15870 33286 0 _0488_
rlabel metal2 16054 30056 16054 30056 0 _0489_
rlabel metal2 16330 30838 16330 30838 0 _0490_
rlabel metal2 15502 32300 15502 32300 0 _0491_
rlabel metal1 16054 33626 16054 33626 0 _0492_
rlabel metal1 14076 32470 14076 32470 0 _0493_
rlabel metal1 15870 32198 15870 32198 0 _0494_
rlabel viali 16361 30668 16361 30668 0 _0495_
rlabel metal1 17572 32402 17572 32402 0 _0496_
rlabel metal2 15318 31280 15318 31280 0 _0497_
rlabel metal1 14628 29818 14628 29818 0 _0498_
rlabel metal1 14628 29138 14628 29138 0 _0499_
rlabel metal2 14306 27200 14306 27200 0 _0500_
rlabel metal1 14168 27574 14168 27574 0 _0501_
rlabel metal1 33028 37094 33028 37094 0 blue
rlabel metal3 1234 13668 1234 13668 0 debug_design_reset
rlabel metal1 14168 37094 14168 37094 0 debug_gpio_ready
rlabel via2 38226 5525 38226 5525 0 design_oeb[0]
rlabel metal1 38778 37094 38778 37094 0 design_oeb[1]
rlabel metal2 25806 1520 25806 1520 0 design_oeb[2]
rlabel metal3 1234 20468 1234 20468 0 design_oeb[3]
rlabel metal3 1234 6868 1234 6868 0 design_oeb[4]
rlabel metal2 32246 1520 32246 1520 0 design_oeb[5]
rlabel metal2 46 1588 46 1588 0 down_key_n
rlabel metal2 6486 1588 6486 1588 0 ext_reset_n
rlabel metal1 7498 23766 7498 23766 0 game.ballDirX
rlabel metal2 9338 27234 9338 27234 0 game.ballDirY
rlabel metal1 6026 24684 6026 24684 0 game.ballX\[0\]
rlabel metal1 10672 25194 10672 25194 0 game.ballX\[1\]
rlabel metal1 7590 23494 7590 23494 0 game.ballX\[2\]
rlabel metal2 12558 21182 12558 21182 0 game.ballX\[3\]
rlabel metal2 2990 20400 2990 20400 0 game.ballX\[4\]
rlabel metal1 5198 17306 5198 17306 0 game.ballX\[5\]
rlabel metal1 8648 18734 8648 18734 0 game.ballX\[6\]
rlabel metal1 7636 16762 7636 16762 0 game.ballX\[7\]
rlabel metal1 5934 21454 5934 21454 0 game.ballX\[8\]
rlabel metal1 7958 26860 7958 26860 0 game.ballY\[0\]
rlabel metal1 8786 27370 8786 27370 0 game.ballY\[1\]
rlabel metal1 5888 28730 5888 28730 0 game.ballY\[2\]
rlabel metal2 3542 28662 3542 28662 0 game.ballY\[3\]
rlabel metal1 8326 30192 8326 30192 0 game.ballY\[4\]
rlabel metal2 6486 31858 6486 31858 0 game.ballY\[5\]
rlabel metal1 9016 32946 9016 32946 0 game.ballY\[6\]
rlabel metal1 10948 32878 10948 32878 0 game.ballY\[7\]
rlabel metal1 23552 21658 23552 21658 0 game.h\[0\]
rlabel metal1 23276 23562 23276 23562 0 game.h\[1\]
rlabel metal2 21022 24820 21022 24820 0 game.h\[2\]
rlabel metal1 23184 24922 23184 24922 0 game.h\[3\]
rlabel metal1 15594 21624 15594 21624 0 game.h\[4\]
rlabel metal1 16606 19890 16606 19890 0 game.h\[5\]
rlabel metal1 21298 20468 21298 20468 0 game.h\[6\]
rlabel metal2 15318 19040 15318 19040 0 game.h\[7\]
rlabel metal1 20148 18666 20148 18666 0 game.h\[8\]
rlabel metal1 14766 19346 14766 19346 0 game.h\[9\]
rlabel via2 14674 31773 14674 31773 0 game.hit
rlabel metal1 13340 24718 13340 24718 0 game.inBallX
rlabel metal2 13570 32241 13570 32241 0 game.inBallY
rlabel metal2 15226 20672 15226 20672 0 game.inPaddle
rlabel metal2 18262 29036 18262 29036 0 game.offset\[0\]
rlabel metal1 20056 31110 20056 31110 0 game.offset\[1\]
rlabel metal2 22034 30804 22034 30804 0 game.offset\[2\]
rlabel metal1 21252 29546 21252 29546 0 game.offset\[3\]
rlabel metal1 21873 27438 21873 27438 0 game.offset\[4\]
rlabel metal2 18446 17442 18446 17442 0 game.paddle\[0\]
rlabel metal1 12834 16116 12834 16116 0 game.paddle\[1\]
rlabel metal2 12834 15640 12834 15640 0 game.paddle\[2\]
rlabel metal1 10028 15470 10028 15470 0 game.paddle\[3\]
rlabel metal1 13110 20366 13110 20366 0 game.paddle\[4\]
rlabel metal2 13570 14178 13570 14178 0 game.paddle\[5\]
rlabel metal2 18814 15878 18814 15878 0 game.paddle\[6\]
rlabel metal1 15548 14042 15548 14042 0 game.paddle\[7\]
rlabel metal1 17020 13498 17020 13498 0 game.paddle\[8\]
rlabel metal1 17940 17782 17940 17782 0 game.v\[0\]
rlabel metal1 18216 26350 18216 26350 0 game.v\[1\]
rlabel metal1 19458 27370 19458 27370 0 game.v\[2\]
rlabel metal1 19550 26316 19550 26316 0 game.v\[3\]
rlabel metal3 15594 20468 15594 20468 0 game.v\[4\]
rlabel metal1 17112 32742 17112 32742 0 game.v\[5\]
rlabel metal1 16238 33354 16238 33354 0 game.v\[6\]
rlabel metal1 16744 32810 16744 32810 0 game.v\[7\]
rlabel metal1 16054 27438 16054 27438 0 game.v\[8\]
rlabel metal1 15134 27948 15134 27948 0 game.v\[9\]
rlabel metal1 20148 37230 20148 37230 0 gpio_ready
rlabel metal2 38686 1520 38686 1520 0 green
rlabel metal2 12926 1520 12926 1520 0 hsync
rlabel metal1 8602 2482 8602 2482 0 net1
rlabel metal1 17687 3094 17687 3094 0 net10
rlabel metal2 19458 37060 19458 37060 0 net11
rlabel metal1 38042 5712 38042 5712 0 net12
rlabel metal1 37950 37230 37950 37230 0 net13
rlabel metal2 25898 2618 25898 2618 0 net14
rlabel metal1 1978 20910 1978 20910 0 net15
rlabel metal1 1702 6970 1702 6970 0 net16
rlabel metal2 32338 2618 32338 2618 0 net17
rlabel metal1 36961 2414 36961 2414 0 net18
rlabel metal1 18009 2482 18009 2482 0 net19
rlabel metal2 6578 7480 6578 7480 0 net2
rlabel metal1 1656 34578 1656 34578 0 net20
rlabel metal2 27186 34612 27186 34612 0 net21
rlabel metal2 1886 27268 1886 27268 0 net22
rlabel metal1 1794 13906 1794 13906 0 net23
rlabel metal1 2530 21012 2530 21012 0 net24
rlabel metal2 1886 18156 1886 18156 0 net25
rlabel metal1 8510 18190 8510 18190 0 net26
rlabel metal1 1794 26350 1794 26350 0 net27
rlabel metal2 8050 24174 8050 24174 0 net28
rlabel metal1 6578 32436 6578 32436 0 net29
rlabel metal1 19872 36754 19872 36754 0 net3
rlabel metal1 2254 31246 2254 31246 0 net30
rlabel metal2 16974 20706 16974 20706 0 net31
rlabel metal1 19734 21998 19734 21998 0 net32
rlabel metal1 18492 17102 18492 17102 0 net33
rlabel metal2 12880 20332 12880 20332 0 net34
rlabel metal1 16054 33014 16054 33014 0 net35
rlabel metal3 15410 31892 15410 31892 0 net36
rlabel metal1 20378 25398 20378 25398 0 net37
rlabel metal1 13754 34034 13754 34034 0 net38
rlabel metal1 2714 31790 2714 31790 0 net39
rlabel metal1 7130 37196 7130 37196 0 net4
rlabel metal2 38318 32793 38318 32793 0 net40
rlabel via2 38318 19125 38318 19125 0 net41
rlabel via2 37766 26333 37766 26333 0 net5
rlabel metal1 19412 2618 19412 2618 0 net6
rlabel metal1 2714 37094 2714 37094 0 net7
rlabel metal2 17066 12478 17066 12478 0 net8
rlabel metal2 32982 34204 32982 34204 0 net9
rlabel metal1 7176 37298 7176 37298 0 new_game_n
rlabel metal3 38234 25908 38234 25908 0 pause_n
rlabel metal3 1234 34068 1234 34068 0 red
rlabel metal1 26910 37094 26910 37094 0 speaker
rlabel metal2 19366 1588 19366 1588 0 up_key_n
rlabel metal3 1234 27268 1234 27268 0 vsync
rlabel metal1 1242 37230 1242 37230 0 wb_clk_i
rlabel metal2 38318 12563 38318 12563 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
