magic
tech sky130A
magscale 1 2
timestamp 1679986744
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37584
<< metal2 >>
rect 662 39200 718 39800
rect 7102 39200 7158 39800
rect 13542 39200 13598 39800
rect 19982 39200 20038 39800
rect 26422 39200 26478 39800
rect 32862 39200 32918 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 6458 200 6514 800
rect 12898 200 12954 800
rect 19338 200 19394 800
rect 25778 200 25834 800
rect 32218 200 32274 800
rect 38658 200 38714 800
<< obsm2 >>
rect 20 39144 606 39200
rect 774 39144 7046 39200
rect 7214 39144 13486 39200
rect 13654 39144 19926 39200
rect 20094 39144 26366 39200
rect 26534 39144 32806 39200
rect 32974 39144 39246 39200
rect 20 856 39356 39144
rect 130 800 6402 856
rect 6570 800 12842 856
rect 13010 800 19282 856
rect 19450 800 25722 856
rect 25890 800 32162 856
rect 32330 800 38602 856
rect 38770 800 39356 856
<< metal3 >>
rect 200 34008 800 34128
rect 39200 32648 39800 32768
rect 200 27208 800 27328
rect 39200 25848 39800 25968
rect 200 20408 800 20528
rect 39200 19048 39800 19168
rect 200 13608 800 13728
rect 39200 12248 39800 12368
rect 200 6808 800 6928
rect 39200 5448 39800 5568
<< obsm3 >>
rect 800 34208 39200 37569
rect 880 33928 39200 34208
rect 800 32848 39200 33928
rect 800 32568 39120 32848
rect 800 27408 39200 32568
rect 880 27128 39200 27408
rect 800 26048 39200 27128
rect 800 25768 39120 26048
rect 800 20608 39200 25768
rect 880 20328 39200 20608
rect 800 19248 39200 20328
rect 800 18968 39120 19248
rect 800 13808 39200 18968
rect 880 13528 39200 13808
rect 800 12448 39200 13528
rect 800 12168 39120 12448
rect 800 7008 39200 12168
rect 880 6728 39200 7008
rect 800 5648 39200 6728
rect 800 5368 39120 5648
rect 800 2143 39200 5368
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 14779 16627 16501 33421
<< labels >>
rlabel metal2 s 32862 39200 32918 39800 6 blue
port 1 nsew signal output
rlabel metal3 s 200 13608 800 13728 6 debug_design_reset
port 2 nsew signal output
rlabel metal2 s 13542 39200 13598 39800 6 debug_gpio_ready
port 3 nsew signal output
rlabel metal3 s 39200 32648 39800 32768 6 debug_oeb[0]
port 4 nsew signal output
rlabel metal3 s 39200 19048 39800 19168 6 debug_oeb[1]
port 5 nsew signal output
rlabel metal3 s 39200 5448 39800 5568 6 design_oeb[0]
port 6 nsew signal output
rlabel metal2 s 39302 39200 39358 39800 6 design_oeb[1]
port 7 nsew signal output
rlabel metal2 s 25778 200 25834 800 6 design_oeb[2]
port 8 nsew signal output
rlabel metal3 s 200 20408 800 20528 6 design_oeb[3]
port 9 nsew signal output
rlabel metal3 s 200 6808 800 6928 6 design_oeb[4]
port 10 nsew signal output
rlabel metal2 s 32218 200 32274 800 6 design_oeb[5]
port 11 nsew signal output
rlabel metal2 s 18 200 74 800 6 down_key_n
port 12 nsew signal input
rlabel metal2 s 6458 200 6514 800 6 ext_reset_n
port 13 nsew signal input
rlabel metal2 s 19982 39200 20038 39800 6 gpio_ready
port 14 nsew signal input
rlabel metal2 s 38658 200 38714 800 6 green
port 15 nsew signal output
rlabel metal2 s 12898 200 12954 800 6 hsync
port 16 nsew signal output
rlabel metal2 s 7102 39200 7158 39800 6 new_game_n
port 17 nsew signal input
rlabel metal3 s 39200 25848 39800 25968 6 pause_n
port 18 nsew signal input
rlabel metal3 s 200 34008 800 34128 6 red
port 19 nsew signal output
rlabel metal2 s 26422 39200 26478 39800 6 speaker
port 20 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 up_key_n
port 21 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 23 nsew ground bidirectional
rlabel metal3 s 200 27208 800 27328 6 vsync
port 24 nsew signal output
rlabel metal2 s 662 39200 718 39800 6 wb_clk_i
port 25 nsew signal input
rlabel metal3 s 39200 12248 39800 12368 6 wb_rst_i
port 26 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2148776
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/solo_squash_caravel/runs/23_03_28_08_55/results/signoff/solo_squash_caravel.magic.gds
string GDS_START 427224
<< end >>

