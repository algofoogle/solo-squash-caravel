// This is the unpowered netlist.
module solo_squash_caravel (blue,
    debug_design_reset,
    debug_gpio_ready,
    down_key_n,
    ext_reset_n,
    gpio_ready,
    green,
    hsync,
    new_game_n,
    pause_n,
    red,
    speaker,
    up_key_n,
    vsync,
    wb_clk_i,
    wb_rst_i,
    debug_oeb,
    design_oeb);
 output blue;
 output debug_design_reset;
 output debug_gpio_ready;
 input down_key_n;
 input ext_reset_n;
 input gpio_ready;
 output green;
 output hsync;
 input new_game_n;
 input pause_n;
 output red;
 output speaker;
 input up_key_n;
 output vsync;
 input wb_clk_i;
 input wb_rst_i;
 output [1:0] debug_oeb;
 output [5:0] design_oeb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire net41;
 wire \game.ballDirX ;
 wire \game.ballDirY ;
 wire \game.ballX[0] ;
 wire \game.ballX[1] ;
 wire \game.ballX[2] ;
 wire \game.ballX[3] ;
 wire \game.ballX[4] ;
 wire \game.ballX[5] ;
 wire \game.ballX[6] ;
 wire \game.ballX[7] ;
 wire \game.ballX[8] ;
 wire \game.ballY[0] ;
 wire \game.ballY[1] ;
 wire \game.ballY[2] ;
 wire \game.ballY[3] ;
 wire \game.ballY[4] ;
 wire \game.ballY[5] ;
 wire \game.ballY[6] ;
 wire \game.ballY[7] ;
 wire \game.h[0] ;
 wire \game.h[1] ;
 wire \game.h[2] ;
 wire \game.h[3] ;
 wire \game.h[4] ;
 wire \game.h[5] ;
 wire \game.h[6] ;
 wire \game.h[7] ;
 wire \game.h[8] ;
 wire \game.h[9] ;
 wire \game.hit ;
 wire \game.inBallX ;
 wire \game.inBallY ;
 wire \game.inPaddle ;
 wire \game.offset[0] ;
 wire \game.offset[1] ;
 wire \game.offset[2] ;
 wire \game.offset[3] ;
 wire \game.offset[4] ;
 wire \game.paddle[0] ;
 wire \game.paddle[1] ;
 wire \game.paddle[2] ;
 wire \game.paddle[3] ;
 wire \game.paddle[4] ;
 wire \game.paddle[5] ;
 wire \game.paddle[6] ;
 wire \game.paddle[7] ;
 wire \game.paddle[8] ;
 wire \game.v[0] ;
 wire \game.v[1] ;
 wire \game.v[2] ;
 wire \game.v[3] ;
 wire \game.v[4] ;
 wire \game.v[5] ;
 wire \game.v[6] ;
 wire \game.v[7] ;
 wire \game.v[8] ;
 wire \game.v[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;

 sky130_fd_sc_hd__and2b_1 _0502_ (.A_N(net8),
    .B(net2),
    .X(_0057_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__clkbuf_2 _0504_ (.A(_0058_),
    .X(_0059_));
 sky130_fd_sc_hd__clkbuf_2 _0505_ (.A(_0059_),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 _0506_ (.A(\game.h[9] ),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_2 _0507_ (.A(\game.h[8] ),
    .X(_0061_));
 sky130_fd_sc_hd__nor3_1 _0508_ (.A(\game.h[5] ),
    .B(\game.h[7] ),
    .C(\game.h[6] ),
    .Y(_0062_));
 sky130_fd_sc_hd__and4bb_1 _0509_ (.A_N(_0060_),
    .B_N(_0061_),
    .C(_0062_),
    .D(\game.inPaddle ),
    .X(_0063_));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(\game.v[4] ),
    .Y(_0064_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0511_ (.A(\game.v[1] ),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_2 _0512_ (.A(_0065_),
    .X(_0066_));
 sky130_fd_sc_hd__or2b_1 _0513_ (.A(\game.v[4] ),
    .B_N(\game.v[3] ),
    .X(_0067_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(_0065_),
    .Y(_0068_));
 sky130_fd_sc_hd__clkinv_2 _0515_ (.A(\game.v[2] ),
    .Y(_0069_));
 sky130_fd_sc_hd__mux2_1 _0516_ (.A0(\game.v[3] ),
    .A1(_0068_),
    .S(_0069_),
    .X(_0070_));
 sky130_fd_sc_hd__o211a_1 _0517_ (.A1(_0064_),
    .A2(_0066_),
    .B1(_0067_),
    .C1(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_2 _0518_ (.A(\game.h[1] ),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_2 _0519_ (.A(\game.h[3] ),
    .X(_0073_));
 sky130_fd_sc_hd__clkbuf_2 _0520_ (.A(\game.h[2] ),
    .X(_0074_));
 sky130_fd_sc_hd__and4_1 _0521_ (.A(_0072_),
    .B(_0073_),
    .C(_0074_),
    .D(\game.h[4] ),
    .X(_0075_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0522_ (.A(_0072_),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_2 _0523_ (.A(\game.h[4] ),
    .X(_0077_));
 sky130_fd_sc_hd__nor4_1 _0524_ (.A(_0076_),
    .B(_0073_),
    .C(_0074_),
    .D(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__buf_2 _0525_ (.A(\game.v[8] ),
    .X(_0079_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0526_ (.A(\game.v[9] ),
    .X(_0080_));
 sky130_fd_sc_hd__a31o_1 _0527_ (.A1(_0079_),
    .A2(\game.v[7] ),
    .A3(\game.v[6] ),
    .B1(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__o21a_1 _0528_ (.A1(\game.h[7] ),
    .A2(\game.h[8] ),
    .B1(\game.h[9] ),
    .X(_0082_));
 sky130_fd_sc_hd__a31o_1 _0529_ (.A1(\game.h[5] ),
    .A2(\game.h[6] ),
    .A3(\game.h[9] ),
    .B1(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__or3_1 _0530_ (.A(\game.v[7] ),
    .B(\game.v[6] ),
    .C(\game.v[5] ),
    .X(_0084_));
 sky130_fd_sc_hd__nor3_1 _0531_ (.A(_0080_),
    .B(_0079_),
    .C(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__or3_1 _0532_ (.A(_0081_),
    .B(_0083_),
    .C(_0085_),
    .X(_0086_));
 sky130_fd_sc_hd__o31a_1 _0533_ (.A1(_0071_),
    .A2(_0075_),
    .A3(_0078_),
    .B1(_0086_),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_2 _0534_ (.A(\game.v[7] ),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_2 _0535_ (.A(\game.v[6] ),
    .X(_0089_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0536_ (.A(\game.v[5] ),
    .X(_0090_));
 sky130_fd_sc_hd__and4_1 _0537_ (.A(_0079_),
    .B(_0088_),
    .C(_0089_),
    .D(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__or3_1 _0538_ (.A(_0080_),
    .B(_0091_),
    .C(_0082_),
    .X(_0092_));
 sky130_fd_sc_hd__o21ba_1 _0539_ (.A1(_0063_),
    .A2(_0087_),
    .B1_N(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_2 _0540_ (.A(_0093_),
    .X(net20));
 sky130_fd_sc_hd__a21oi_2 _0541_ (.A1(\game.inBallY ),
    .A2(\game.inBallX ),
    .B1(_0086_),
    .Y(_0094_));
 sky130_fd_sc_hd__nor2_2 _0542_ (.A(_0092_),
    .B(_0094_),
    .Y(net18));
 sky130_fd_sc_hd__clkbuf_2 _0543_ (.A(\game.v[2] ),
    .X(_0095_));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(\game.v[9] ),
    .Y(_0096_));
 sky130_fd_sc_hd__nand2_1 _0545_ (.A(_0096_),
    .B(_0091_),
    .Y(_0097_));
 sky130_fd_sc_hd__or4_1 _0546_ (.A(_0095_),
    .B(_0068_),
    .C(_0067_),
    .D(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0547_ (.A(_0098_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 _0548_ (.A(\game.h[5] ),
    .X(_0099_));
 sky130_fd_sc_hd__and3_1 _0549_ (.A(_0099_),
    .B(_0077_),
    .C(\game.h[6] ),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _0550_ (.A(\game.h[7] ),
    .B(_0060_),
    .Y(_0101_));
 sky130_fd_sc_hd__or3_1 _0551_ (.A(_0099_),
    .B(_0077_),
    .C(\game.h[6] ),
    .X(_0102_));
 sky130_fd_sc_hd__or4b_1 _0552_ (.A(_0061_),
    .B(_0100_),
    .C(_0101_),
    .D_N(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_1 _0553_ (.A(_0103_),
    .X(net19));
 sky130_fd_sc_hd__buf_2 _0554_ (.A(\game.v[3] ),
    .X(_0104_));
 sky130_fd_sc_hd__inv_2 _0555_ (.A(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2_1 _0556_ (.A(_0105_),
    .B(\game.offset[4] ),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(\game.offset[3] ),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _0558_ (.A(\game.v[0] ),
    .Y(_0108_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0559_ (.A(\game.offset[2] ),
    .X(_0109_));
 sky130_fd_sc_hd__or2b_1 _0560_ (.A(_0109_),
    .B_N(_0065_),
    .X(_0110_));
 sky130_fd_sc_hd__and2b_1 _0561_ (.A_N(_0065_),
    .B(_0109_),
    .X(_0111_));
 sky130_fd_sc_hd__a31o_1 _0562_ (.A1(_0108_),
    .A2(\game.offset[1] ),
    .A3(_0110_),
    .B1(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__a21oi_1 _0563_ (.A1(_0069_),
    .A2(\game.offset[3] ),
    .B1(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__a21o_1 _0564_ (.A1(_0095_),
    .A2(_0107_),
    .B1(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__nor2_1 _0565_ (.A(_0105_),
    .B(\game.offset[4] ),
    .Y(_0115_));
 sky130_fd_sc_hd__a21oi_1 _0566_ (.A1(_0106_),
    .A2(_0114_),
    .B1(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__or2b_1 _0567_ (.A(_0073_),
    .B_N(\game.offset[4] ),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _0568_ (.A(_0107_),
    .B(\game.h[2] ),
    .X(_0118_));
 sky130_fd_sc_hd__or2b_1 _0569_ (.A(_0072_),
    .B_N(\game.offset[2] ),
    .X(_0119_));
 sky130_fd_sc_hd__or2b_1 _0570_ (.A(\game.h[0] ),
    .B_N(\game.offset[1] ),
    .X(_0120_));
 sky130_fd_sc_hd__and2b_1 _0571_ (.A_N(\game.offset[2] ),
    .B(_0072_),
    .X(_0121_));
 sky130_fd_sc_hd__a21o_1 _0572_ (.A1(_0119_),
    .A2(_0120_),
    .B1(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__and2_1 _0573_ (.A(_0107_),
    .B(\game.h[2] ),
    .X(_0123_));
 sky130_fd_sc_hd__a21o_1 _0574_ (.A1(_0118_),
    .A2(_0122_),
    .B1(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__and2b_1 _0575_ (.A_N(\game.offset[4] ),
    .B(_0073_),
    .X(_0125_));
 sky130_fd_sc_hd__a21oi_1 _0576_ (.A1(_0117_),
    .A2(_0124_),
    .B1(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__clkbuf_2 _0577_ (.A(\game.v[4] ),
    .X(_0127_));
 sky130_fd_sc_hd__xnor2_1 _0578_ (.A(_0127_),
    .B(_0077_),
    .Y(_0128_));
 sky130_fd_sc_hd__xnor2_1 _0579_ (.A(_0126_),
    .B(_0128_),
    .Y(_0129_));
 sky130_fd_sc_hd__xnor2_1 _0580_ (.A(_0116_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__clkbuf_2 _0581_ (.A(\game.v[0] ),
    .X(_0131_));
 sky130_fd_sc_hd__xnor2_1 _0582_ (.A(_0131_),
    .B(\game.offset[1] ),
    .Y(_0132_));
 sky130_fd_sc_hd__xnor2_1 _0583_ (.A(_0131_),
    .B(\game.h[0] ),
    .Y(_0133_));
 sky130_fd_sc_hd__o21a_1 _0584_ (.A1(_0130_),
    .A2(_0132_),
    .B1(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__xnor2_1 _0585_ (.A(\game.v[2] ),
    .B(_0074_),
    .Y(_0135_));
 sky130_fd_sc_hd__xnor2_1 _0586_ (.A(_0112_),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__xnor2_1 _0587_ (.A(_0124_),
    .B(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__xor2_1 _0588_ (.A(\game.v[3] ),
    .B(\game.h[3] ),
    .X(_0138_));
 sky130_fd_sc_hd__xnor2_1 _0589_ (.A(_0122_),
    .B(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__xnor2_1 _0590_ (.A(_0114_),
    .B(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__xnor2_1 _0591_ (.A(_0137_),
    .B(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__a21oi_1 _0592_ (.A1(_0133_),
    .A2(_0141_),
    .B1(_0130_),
    .Y(_0142_));
 sky130_fd_sc_hd__a21bo_1 _0593_ (.A1(_0130_),
    .A2(_0141_),
    .B1_N(_0094_),
    .X(_0143_));
 sky130_fd_sc_hd__nor4_1 _0594_ (.A(net20),
    .B(_0134_),
    .C(_0142_),
    .D(_0143_),
    .Y(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0595_ (.A(\game.ballY[5] ),
    .X(_0144_));
 sky130_fd_sc_hd__nor2_1 _0596_ (.A(\game.ballY[4] ),
    .B(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0597_ (.A(\game.ballY[6] ),
    .X(_0146_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0598_ (.A(\game.ballY[7] ),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_1 _0599_ (.A(_0146_),
    .B(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__clkbuf_2 _0600_ (.A(\game.ballY[3] ),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _0601_ (.A(_0149_),
    .B(\game.ballY[4] ),
    .X(_0150_));
 sky130_fd_sc_hd__o211a_1 _0602_ (.A1(_0144_),
    .A2(_0150_),
    .B1(_0147_),
    .C1(_0146_),
    .X(_0151_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0603_ (.A(\game.ballX[6] ),
    .X(_0152_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0604_ (.A(\game.ballX[7] ),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_2 _0605_ (.A(\game.ballX[4] ),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_2 _0606_ (.A(\game.ballX[5] ),
    .X(_0155_));
 sky130_fd_sc_hd__o21a_1 _0607_ (.A1(\game.ballX[3] ),
    .A2(_0154_),
    .B1(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__o31a_1 _0608_ (.A1(_0152_),
    .A2(_0153_),
    .A3(_0156_),
    .B1(\game.ballX[8] ),
    .X(_0157_));
 sky130_fd_sc_hd__a211o_1 _0609_ (.A1(_0145_),
    .A2(_0148_),
    .B1(_0151_),
    .C1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0610_ (.A(_0089_),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _0611_ (.A1(_0090_),
    .A2(\game.hit ),
    .B1(_0158_),
    .B2(_0159_),
    .X(net21));
 sky130_fd_sc_hd__and4_1 _0612_ (.A(\game.h[1] ),
    .B(\game.h[0] ),
    .C(\game.h[3] ),
    .D(\game.h[2] ),
    .X(_0160_));
 sky130_fd_sc_hd__and2_1 _0613_ (.A(\game.h[4] ),
    .B(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__nand4_2 _0614_ (.A(_0060_),
    .B(_0061_),
    .C(_0062_),
    .D(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__or4bb_1 _0615_ (.A(\game.v[1] ),
    .B(\game.v[0] ),
    .C_N(\game.v[3] ),
    .D_N(\game.v[2] ),
    .X(_0163_));
 sky130_fd_sc_hd__or4b_1 _0616_ (.A(\game.v[8] ),
    .B(\game.v[5] ),
    .C(\game.v[4] ),
    .D_N(\game.v[9] ),
    .X(_0164_));
 sky130_fd_sc_hd__nor4_1 _0617_ (.A(\game.v[7] ),
    .B(\game.v[6] ),
    .C(_0163_),
    .D(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand2_1 _0618_ (.A(net5),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__nor2_2 _0619_ (.A(_0162_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__clkbuf_2 _0620_ (.A(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__and4_1 _0621_ (.A(\game.h[9] ),
    .B(\game.h[8] ),
    .C(_0062_),
    .D(_0161_),
    .X(_0169_));
 sky130_fd_sc_hd__or4_1 _0622_ (.A(_0096_),
    .B(_0069_),
    .C(_0065_),
    .D(\game.v[0] ),
    .X(_0170_));
 sky130_fd_sc_hd__nor4_1 _0623_ (.A(\game.v[8] ),
    .B(_0084_),
    .C(_0067_),
    .D(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__and3_1 _0624_ (.A(net5),
    .B(_0169_),
    .C(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__buf_2 _0625_ (.A(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__nand2_1 _0626_ (.A(\game.offset[0] ),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__clkbuf_2 _0627_ (.A(_0057_),
    .X(_0175_));
 sky130_fd_sc_hd__buf_2 _0628_ (.A(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__o211a_1 _0629_ (.A1(\game.offset[0] ),
    .A2(_0168_),
    .B1(_0174_),
    .C1(_0176_),
    .X(_0000_));
 sky130_fd_sc_hd__and3_1 _0630_ (.A(\game.offset[1] ),
    .B(\game.offset[0] ),
    .C(_0167_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_2 _0631_ (.A(_0057_),
    .X(_0178_));
 sky130_fd_sc_hd__a21o_1 _0632_ (.A1(\game.offset[0] ),
    .A2(_0167_),
    .B1(\game.offset[1] ),
    .X(_0179_));
 sky130_fd_sc_hd__and3b_1 _0633_ (.A_N(_0177_),
    .B(_0178_),
    .C(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _0634_ (.A(_0180_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _0635_ (.A(_0109_),
    .B(_0177_),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _0636_ (.A(_0109_),
    .B(_0177_),
    .Y(_0182_));
 sky130_fd_sc_hd__and3_1 _0637_ (.A(_0175_),
    .B(_0181_),
    .C(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _0638_ (.A(_0183_),
    .X(_0002_));
 sky130_fd_sc_hd__and3_1 _0639_ (.A(\game.offset[3] ),
    .B(_0109_),
    .C(_0177_),
    .X(_0184_));
 sky130_fd_sc_hd__a21o_1 _0640_ (.A1(_0109_),
    .A2(_0177_),
    .B1(\game.offset[3] ),
    .X(_0185_));
 sky130_fd_sc_hd__and3b_1 _0641_ (.A_N(_0184_),
    .B(_0178_),
    .C(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0642_ (.A(_0186_),
    .X(_0003_));
 sky130_fd_sc_hd__xnor2_1 _0643_ (.A(\game.offset[4] ),
    .B(_0184_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _0644_ (.A(net24),
    .B(_0187_),
    .Y(_0004_));
 sky130_fd_sc_hd__clkbuf_2 _0645_ (.A(net4),
    .X(_0188_));
 sky130_fd_sc_hd__or4_1 _0646_ (.A(_0096_),
    .B(\game.v[8] ),
    .C(_0084_),
    .D(_0067_),
    .X(_0189_));
 sky130_fd_sc_hd__and4bb_1 _0647_ (.A_N(_0066_),
    .B_N(_0189_),
    .C(_0108_),
    .D(_0095_),
    .X(_0190_));
 sky130_fd_sc_hd__and3_1 _0648_ (.A(net5),
    .B(_0169_),
    .C(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_2 _0649_ (.A(\game.paddle[8] ),
    .X(_0192_));
 sky130_fd_sc_hd__a21oi_1 _0650_ (.A1(\game.paddle[7] ),
    .A2(_0192_),
    .B1(net1),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _0651_ (.A(net6),
    .Y(_0194_));
 sky130_fd_sc_hd__o41a_1 _0652_ (.A1(\game.paddle[5] ),
    .A2(\game.paddle[6] ),
    .A3(\game.paddle[7] ),
    .A4(\game.paddle[8] ),
    .B1(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__or2_1 _0653_ (.A(_0193_),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__and2_1 _0654_ (.A(_0191_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _0655_ (.A(_0188_),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__and3_1 _0656_ (.A(\game.paddle[0] ),
    .B(_0178_),
    .C(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _0657_ (.A(_0199_),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_2 _0658_ (.A(_0057_),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_1 _0659_ (.A(_0173_),
    .B(_0196_),
    .Y(_0201_));
 sky130_fd_sc_hd__and2_1 _0660_ (.A(net4),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_2 _0661_ (.A(\game.paddle[1] ),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0662_ (.A0(_0197_),
    .A1(_0202_),
    .S(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__and2_1 _0663_ (.A(_0200_),
    .B(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _0664_ (.A(_0205_),
    .X(_0006_));
 sky130_fd_sc_hd__clkbuf_2 _0665_ (.A(\game.paddle[2] ),
    .X(_0206_));
 sky130_fd_sc_hd__or2_2 _0666_ (.A(_0162_),
    .B(_0166_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_2 _0667_ (.A(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__a21o_1 _0668_ (.A1(\game.paddle[7] ),
    .A2(_0192_),
    .B1(net1),
    .X(_0209_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0669_ (.A(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _0670_ (.A(_0209_),
    .B(_0195_),
    .Y(_0211_));
 sky130_fd_sc_hd__xor2_1 _0671_ (.A(\game.paddle[1] ),
    .B(_0206_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _0672_ (.A0(_0210_),
    .A1(_0211_),
    .S(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__or2_1 _0673_ (.A(_0208_),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__o21a_1 _0674_ (.A1(_0206_),
    .A2(_0197_),
    .B1(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _0675_ (.A(_0175_),
    .B(_0198_),
    .C(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _0676_ (.A(_0216_),
    .X(_0007_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0677_ (.A(\game.paddle[3] ),
    .X(_0217_));
 sky130_fd_sc_hd__o21ai_1 _0678_ (.A1(_0203_),
    .A2(_0206_),
    .B1(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__or3_1 _0679_ (.A(\game.paddle[1] ),
    .B(\game.paddle[2] ),
    .C(_0217_),
    .X(_0219_));
 sky130_fd_sc_hd__and2_1 _0680_ (.A(_0218_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__a31o_1 _0681_ (.A1(_0203_),
    .A2(_0206_),
    .A3(_0217_),
    .B1(_0210_),
    .X(_0221_));
 sky130_fd_sc_hd__a21oi_1 _0682_ (.A1(_0203_),
    .A2(_0206_),
    .B1(_0217_),
    .Y(_0222_));
 sky130_fd_sc_hd__o22a_1 _0683_ (.A1(_0211_),
    .A2(_0220_),
    .B1(_0221_),
    .B2(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_2 _0684_ (.A(_0208_),
    .X(_0224_));
 sky130_fd_sc_hd__o2bb2a_1 _0685_ (.A1_N(_0217_),
    .A2_N(_0202_),
    .B1(_0223_),
    .B2(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__nor2_1 _0686_ (.A(net23),
    .B(_0225_),
    .Y(_0008_));
 sky130_fd_sc_hd__a21bo_1 _0687_ (.A1(_0210_),
    .A2(_0219_),
    .B1_N(_0221_),
    .X(_0226_));
 sky130_fd_sc_hd__xor2_1 _0688_ (.A(\game.paddle[4] ),
    .B(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _0689_ (.A(_0201_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__a21oi_1 _0690_ (.A1(\game.paddle[4] ),
    .A2(_0202_),
    .B1(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__nor2_1 _0691_ (.A(net23),
    .B(_0229_),
    .Y(_0009_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0692_ (.A(\game.paddle[5] ),
    .X(_0230_));
 sky130_fd_sc_hd__or3_1 _0693_ (.A(\game.paddle[4] ),
    .B(_0230_),
    .C(_0219_),
    .X(_0231_));
 sky130_fd_sc_hd__o21ai_1 _0694_ (.A1(\game.paddle[4] ),
    .A2(_0219_),
    .B1(_0230_),
    .Y(_0232_));
 sky130_fd_sc_hd__and2_1 _0695_ (.A(_0231_),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__and4_1 _0696_ (.A(\game.paddle[1] ),
    .B(\game.paddle[2] ),
    .C(\game.paddle[3] ),
    .D(\game.paddle[4] ),
    .X(_0234_));
 sky130_fd_sc_hd__and2_1 _0697_ (.A(\game.paddle[5] ),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _0698_ (.A(_0209_),
    .B(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_1 _0699_ (.A(_0230_),
    .B(_0234_),
    .Y(_0237_));
 sky130_fd_sc_hd__o22a_1 _0700_ (.A1(_0211_),
    .A2(_0233_),
    .B1(_0236_),
    .B2(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__o2bb2a_1 _0701_ (.A1_N(_0230_),
    .A2_N(_0202_),
    .B1(_0238_),
    .B2(_0224_),
    .X(_0239_));
 sky130_fd_sc_hd__nor2_1 _0702_ (.A(net23),
    .B(_0239_),
    .Y(_0010_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0703_ (.A(\game.paddle[6] ),
    .X(_0240_));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(_0236_),
    .Y(_0241_));
 sky130_fd_sc_hd__a211o_1 _0705_ (.A1(_0210_),
    .A2(_0231_),
    .B1(_0241_),
    .C1(_0201_),
    .X(_0242_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(\game.paddle[6] ),
    .Y(_0243_));
 sky130_fd_sc_hd__a21bo_1 _0707_ (.A1(_0243_),
    .A2(_0198_),
    .B1_N(_0242_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_2 _0708_ (.A(_0057_),
    .X(_0245_));
 sky130_fd_sc_hd__o211ai_1 _0709_ (.A1(_0240_),
    .A2(_0242_),
    .B1(_0244_),
    .C1(_0245_),
    .Y(_0011_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0710_ (.A(\game.paddle[7] ),
    .X(_0246_));
 sky130_fd_sc_hd__o2bb2a_1 _0711_ (.A1_N(_0240_),
    .A2_N(_0235_),
    .B1(_0231_),
    .B2(_0193_),
    .X(_0247_));
 sky130_fd_sc_hd__a211oi_1 _0712_ (.A1(_0240_),
    .A2(_0210_),
    .B1(_0201_),
    .C1(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _0713_ (.A(_0246_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__o2111a_1 _0714_ (.A1(_0246_),
    .A2(_0248_),
    .B1(_0249_),
    .C1(_0245_),
    .D1(_0198_),
    .X(_0012_));
 sky130_fd_sc_hd__nor3_1 _0715_ (.A(_0240_),
    .B(_0246_),
    .C(_0231_),
    .Y(_0250_));
 sky130_fd_sc_hd__a31o_1 _0716_ (.A1(_0240_),
    .A2(_0246_),
    .A3(_0235_),
    .B1(_0210_),
    .X(_0251_));
 sky130_fd_sc_hd__o21a_1 _0717_ (.A1(_0193_),
    .A2(_0250_),
    .B1(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__a22oi_1 _0718_ (.A1(_0192_),
    .A2(_0198_),
    .B1(_0252_),
    .B2(_0197_),
    .Y(_0253_));
 sky130_fd_sc_hd__a31o_1 _0719_ (.A1(_0192_),
    .A2(_0197_),
    .A3(_0252_),
    .B1(_0059_),
    .X(_0254_));
 sky130_fd_sc_hd__nor2_1 _0720_ (.A(_0253_),
    .B(_0254_),
    .Y(_0013_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0721_ (.A(\game.ballY[0] ),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _0722_ (.A(net4),
    .B(_0207_),
    .Y(_0256_));
 sky130_fd_sc_hd__clkbuf_2 _0723_ (.A(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _0724_ (.A(_0255_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__o211a_1 _0725_ (.A1(_0255_),
    .A2(_0168_),
    .B1(_0258_),
    .C1(_0176_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _0726_ (.A(net4),
    .B(_0207_),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_2 _0727_ (.A(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_1 _0728_ (.A(\game.ballY[1] ),
    .B(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_1 _0729_ (.A(\game.ballDirY ),
    .B(\game.ballY[1] ),
    .Y(_0262_));
 sky130_fd_sc_hd__or2_1 _0730_ (.A(\game.ballDirY ),
    .B(\game.ballY[1] ),
    .X(_0263_));
 sky130_fd_sc_hd__a21oi_1 _0731_ (.A1(_0262_),
    .A2(_0263_),
    .B1(_0255_),
    .Y(_0264_));
 sky130_fd_sc_hd__and3_1 _0732_ (.A(_0255_),
    .B(_0262_),
    .C(_0263_),
    .X(_0265_));
 sky130_fd_sc_hd__or3_1 _0733_ (.A(_0208_),
    .B(_0264_),
    .C(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__clkbuf_2 _0734_ (.A(_0059_),
    .X(_0267_));
 sky130_fd_sc_hd__a21oi_1 _0735_ (.A1(_0261_),
    .A2(_0266_),
    .B1(_0267_),
    .Y(_0015_));
 sky130_fd_sc_hd__clkbuf_2 _0736_ (.A(_0059_),
    .X(_0268_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0737_ (.A(\game.ballDirY ),
    .X(_0269_));
 sky130_fd_sc_hd__or2b_1 _0738_ (.A(\game.ballY[2] ),
    .B_N(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__or2b_1 _0739_ (.A(\game.ballDirY ),
    .B_N(\game.ballY[2] ),
    .X(_0271_));
 sky130_fd_sc_hd__a21bo_1 _0740_ (.A1(\game.ballY[0] ),
    .A2(_0263_),
    .B1_N(_0262_),
    .X(_0272_));
 sky130_fd_sc_hd__a21o_1 _0741_ (.A1(_0270_),
    .A2(_0271_),
    .B1(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__nand3_1 _0742_ (.A(_0270_),
    .B(_0271_),
    .C(_0272_),
    .Y(_0274_));
 sky130_fd_sc_hd__and3_1 _0743_ (.A(_0168_),
    .B(_0273_),
    .C(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__a21oi_1 _0744_ (.A1(\game.ballY[2] ),
    .A2(_0260_),
    .B1(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2_1 _0745_ (.A(_0268_),
    .B(_0276_),
    .Y(_0016_));
 sky130_fd_sc_hd__or2b_1 _0746_ (.A(\game.ballY[3] ),
    .B_N(\game.ballDirY ),
    .X(_0277_));
 sky130_fd_sc_hd__or2b_1 _0747_ (.A(_0269_),
    .B_N(_0149_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_1 _0748_ (.A(_0277_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__a21oi_1 _0749_ (.A1(_0271_),
    .A2(_0274_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__and3_1 _0750_ (.A(_0271_),
    .B(_0274_),
    .C(_0279_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _0751_ (.A(_0280_),
    .B(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__o2bb2a_1 _0752_ (.A1_N(_0149_),
    .A2_N(_0260_),
    .B1(_0282_),
    .B2(_0224_),
    .X(_0283_));
 sky130_fd_sc_hd__nor2_1 _0753_ (.A(_0268_),
    .B(_0283_),
    .Y(_0017_));
 sky130_fd_sc_hd__o21ba_1 _0754_ (.A1(\game.ballY[2] ),
    .A2(\game.ballY[3] ),
    .B1_N(_0269_),
    .X(_0284_));
 sky130_fd_sc_hd__a41o_1 _0755_ (.A1(_0270_),
    .A2(_0271_),
    .A3(_0272_),
    .A4(_0277_),
    .B1(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__xnor2_1 _0756_ (.A(_0269_),
    .B(\game.ballY[4] ),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_1 _0757_ (.A(_0285_),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__o21a_1 _0758_ (.A1(_0285_),
    .A2(_0286_),
    .B1(_0173_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(\game.ballY[4] ),
    .Y(_0289_));
 sky130_fd_sc_hd__o2bb2a_1 _0760_ (.A1_N(_0287_),
    .A2_N(_0288_),
    .B1(_0289_),
    .B2(_0257_),
    .X(_0290_));
 sky130_fd_sc_hd__nor2_1 _0761_ (.A(_0268_),
    .B(_0290_),
    .Y(_0018_));
 sky130_fd_sc_hd__nor2_1 _0762_ (.A(_0144_),
    .B(_0257_),
    .Y(_0291_));
 sky130_fd_sc_hd__clkbuf_2 _0763_ (.A(_0269_),
    .X(_0292_));
 sky130_fd_sc_hd__o21ai_1 _0764_ (.A1(_0292_),
    .A2(_0289_),
    .B1(_0287_),
    .Y(_0293_));
 sky130_fd_sc_hd__xor2_1 _0765_ (.A(\game.ballDirY ),
    .B(\game.ballY[5] ),
    .X(_0294_));
 sky130_fd_sc_hd__o21ai_1 _0766_ (.A1(_0293_),
    .A2(_0294_),
    .B1(_0173_),
    .Y(_0295_));
 sky130_fd_sc_hd__a21oi_1 _0767_ (.A1(_0293_),
    .A2(_0294_),
    .B1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__o21ai_1 _0768_ (.A1(_0291_),
    .A2(_0296_),
    .B1(_0176_),
    .Y(_0019_));
 sky130_fd_sc_hd__xnor2_1 _0769_ (.A(_0292_),
    .B(_0146_),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(_0294_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _0771_ (.A(_0269_),
    .B(_0145_),
    .Y(_0299_));
 sky130_fd_sc_hd__a31o_1 _0772_ (.A1(_0285_),
    .A2(_0286_),
    .A3(_0298_),
    .B1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2_1 _0773_ (.A(_0297_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__or2_1 _0774_ (.A(_0297_),
    .B(_0300_),
    .X(_0302_));
 sky130_fd_sc_hd__and3_1 _0775_ (.A(_0188_),
    .B(_0146_),
    .C(_0208_),
    .X(_0303_));
 sky130_fd_sc_hd__a31o_1 _0776_ (.A1(_0168_),
    .A2(_0301_),
    .A3(_0302_),
    .B1(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__and2_1 _0777_ (.A(_0200_),
    .B(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _0778_ (.A(_0305_),
    .X(_0020_));
 sky130_fd_sc_hd__or2b_1 _0779_ (.A(_0292_),
    .B_N(_0146_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _0780_ (.A(_0292_),
    .B(_0147_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_1 _0781_ (.A(_0292_),
    .B(_0147_),
    .Y(_0308_));
 sky130_fd_sc_hd__a22o_1 _0782_ (.A1(_0306_),
    .A2(_0301_),
    .B1(_0307_),
    .B2(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__nand4_1 _0783_ (.A(_0306_),
    .B(_0301_),
    .C(_0307_),
    .D(_0308_),
    .Y(_0310_));
 sky130_fd_sc_hd__and3_1 _0784_ (.A(_0188_),
    .B(_0147_),
    .C(_0207_),
    .X(_0311_));
 sky130_fd_sc_hd__a31o_1 _0785_ (.A1(_0167_),
    .A2(_0309_),
    .A3(_0310_),
    .B1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__and2_1 _0786_ (.A(_0200_),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _0787_ (.A(_0313_),
    .X(_0021_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0788_ (.A(\game.ballX[0] ),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _0789_ (.A(_0314_),
    .B(_0257_),
    .Y(_0315_));
 sky130_fd_sc_hd__o211a_1 _0790_ (.A1(_0314_),
    .A2(_0168_),
    .B1(_0315_),
    .C1(_0176_),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _0791_ (.A(\game.ballX[1] ),
    .B(_0260_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _0792_ (.A(\game.ballDirX ),
    .B(\game.ballX[1] ),
    .Y(_0317_));
 sky130_fd_sc_hd__or2_1 _0793_ (.A(\game.ballDirX ),
    .B(\game.ballX[1] ),
    .X(_0318_));
 sky130_fd_sc_hd__a21oi_1 _0794_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0314_),
    .Y(_0319_));
 sky130_fd_sc_hd__and3_1 _0795_ (.A(_0314_),
    .B(_0317_),
    .C(_0318_),
    .X(_0320_));
 sky130_fd_sc_hd__or3_1 _0796_ (.A(_0208_),
    .B(_0319_),
    .C(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__a21oi_1 _0797_ (.A1(_0316_),
    .A2(_0321_),
    .B1(_0267_),
    .Y(_0023_));
 sky130_fd_sc_hd__clkbuf_2 _0798_ (.A(\game.ballDirX ),
    .X(_0322_));
 sky130_fd_sc_hd__or2b_1 _0799_ (.A(\game.ballX[2] ),
    .B_N(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_2 _0800_ (.A(_0322_),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_2 _0801_ (.A(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or2b_1 _0802_ (.A(_0325_),
    .B_N(\game.ballX[2] ),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _0803_ (.A(_0323_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21bo_1 _0804_ (.A1(\game.ballX[0] ),
    .A2(_0318_),
    .B1_N(_0317_),
    .X(_0328_));
 sky130_fd_sc_hd__xor2_1 _0805_ (.A(_0327_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__o2bb2a_1 _0806_ (.A1_N(\game.ballX[2] ),
    .A2_N(_0260_),
    .B1(_0329_),
    .B2(_0224_),
    .X(_0330_));
 sky130_fd_sc_hd__nor2_1 _0807_ (.A(_0268_),
    .B(_0330_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(\game.ballX[3] ),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2_1 _0809_ (.A(_0322_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__or2_1 _0810_ (.A(_0325_),
    .B(_0331_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _0811_ (.A(_0332_),
    .B(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__and2b_1 _0812_ (.A_N(_0322_),
    .B(\game.ballX[2] ),
    .X(_0335_));
 sky130_fd_sc_hd__a21oi_1 _0813_ (.A1(_0323_),
    .A2(_0328_),
    .B1(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__xnor2_1 _0814_ (.A(_0334_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__o22a_1 _0815_ (.A1(_0331_),
    .A2(_0257_),
    .B1(_0337_),
    .B2(_0224_),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_1 _0816_ (.A(_0268_),
    .B(_0338_),
    .Y(_0025_));
 sky130_fd_sc_hd__xnor2_1 _0817_ (.A(_0324_),
    .B(\game.ballX[4] ),
    .Y(_0339_));
 sky130_fd_sc_hd__nor2_1 _0818_ (.A(_0322_),
    .B(_0331_),
    .Y(_0340_));
 sky130_fd_sc_hd__a311o_1 _0819_ (.A1(_0323_),
    .A2(_0328_),
    .A3(_0332_),
    .B1(_0340_),
    .C1(_0335_),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _0820_ (.A(_0339_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__o21a_1 _0821_ (.A1(_0339_),
    .A2(_0341_),
    .B1(_0173_),
    .X(_0343_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(\game.ballX[4] ),
    .Y(_0344_));
 sky130_fd_sc_hd__o2bb2a_1 _0823_ (.A1_N(_0342_),
    .A2_N(_0343_),
    .B1(_0344_),
    .B2(_0257_),
    .X(_0345_));
 sky130_fd_sc_hd__nor2_1 _0824_ (.A(_0268_),
    .B(_0345_),
    .Y(_0026_));
 sky130_fd_sc_hd__xor2_1 _0825_ (.A(_0322_),
    .B(\game.ballX[5] ),
    .X(_0346_));
 sky130_fd_sc_hd__o21ai_1 _0826_ (.A1(_0325_),
    .A2(_0344_),
    .B1(_0342_),
    .Y(_0347_));
 sky130_fd_sc_hd__and2_1 _0827_ (.A(_0346_),
    .B(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__o21ai_1 _0828_ (.A1(_0346_),
    .A2(_0347_),
    .B1(_0173_),
    .Y(_0349_));
 sky130_fd_sc_hd__o22a_1 _0829_ (.A1(_0155_),
    .A2(_0256_),
    .B1(_0348_),
    .B2(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _0830_ (.A(_0059_),
    .B(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0831_ (.A(_0351_),
    .X(_0027_));
 sky130_fd_sc_hd__and3_1 _0832_ (.A(_0188_),
    .B(_0152_),
    .C(_0224_),
    .X(_0352_));
 sky130_fd_sc_hd__xnor2_1 _0833_ (.A(_0324_),
    .B(\game.ballX[6] ),
    .Y(_0353_));
 sky130_fd_sc_hd__clkinv_2 _0834_ (.A(_0346_),
    .Y(_0354_));
 sky130_fd_sc_hd__and3_1 _0835_ (.A(_0339_),
    .B(_0341_),
    .C(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__o21ba_1 _0836_ (.A1(_0154_),
    .A2(_0155_),
    .B1_N(_0324_),
    .X(_0356_));
 sky130_fd_sc_hd__or3_1 _0837_ (.A(_0353_),
    .B(_0355_),
    .C(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__o21ai_1 _0838_ (.A1(_0355_),
    .A2(_0356_),
    .B1(_0353_),
    .Y(_0358_));
 sky130_fd_sc_hd__and3_1 _0839_ (.A(_0168_),
    .B(_0357_),
    .C(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__o21a_1 _0840_ (.A1(_0352_),
    .A2(_0359_),
    .B1(_0176_),
    .X(_0028_));
 sky130_fd_sc_hd__xnor2_1 _0841_ (.A(_0324_),
    .B(\game.ballX[7] ),
    .Y(_0360_));
 sky130_fd_sc_hd__or2b_1 _0842_ (.A(_0325_),
    .B_N(_0152_),
    .X(_0361_));
 sky130_fd_sc_hd__nand3b_1 _0843_ (.A_N(_0360_),
    .B(_0358_),
    .C(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__a21bo_1 _0844_ (.A1(_0361_),
    .A2(_0358_),
    .B1_N(_0360_),
    .X(_0363_));
 sky130_fd_sc_hd__and3_1 _0845_ (.A(_0188_),
    .B(_0153_),
    .C(_0207_),
    .X(_0364_));
 sky130_fd_sc_hd__a31o_1 _0846_ (.A1(_0167_),
    .A2(_0362_),
    .A3(_0363_),
    .B1(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__and2_1 _0847_ (.A(_0200_),
    .B(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0366_),
    .X(_0029_));
 sky130_fd_sc_hd__nand2_1 _0849_ (.A(\game.ballX[8] ),
    .B(_0260_),
    .Y(_0367_));
 sky130_fd_sc_hd__and3_1 _0850_ (.A(_0353_),
    .B(_0355_),
    .C(_0360_),
    .X(_0368_));
 sky130_fd_sc_hd__o21ba_1 _0851_ (.A1(_0152_),
    .A2(_0153_),
    .B1_N(_0324_),
    .X(_0369_));
 sky130_fd_sc_hd__xnor2_1 _0852_ (.A(_0325_),
    .B(\game.ballX[8] ),
    .Y(_0370_));
 sky130_fd_sc_hd__o31a_1 _0853_ (.A1(_0356_),
    .A2(_0368_),
    .A3(_0369_),
    .B1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__or4_1 _0854_ (.A(_0356_),
    .B(_0368_),
    .C(_0369_),
    .D(_0370_),
    .X(_0372_));
 sky130_fd_sc_hd__or3b_1 _0855_ (.A(_0371_),
    .B(_0208_),
    .C_N(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__a21oi_1 _0856_ (.A1(_0367_),
    .A2(_0373_),
    .B1(_0267_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(_0217_),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _0858_ (.A(\game.v[5] ),
    .Y(_0375_));
 sky130_fd_sc_hd__o22a_1 _0859_ (.A1(_0069_),
    .A2(\game.paddle[2] ),
    .B1(_0230_),
    .B2(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__o221ai_1 _0860_ (.A1(_0068_),
    .A2(_0203_),
    .B1(_0374_),
    .B2(_0104_),
    .C1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__xor2_1 _0861_ (.A(\game.v[0] ),
    .B(\game.paddle[0] ),
    .X(_0378_));
 sky130_fd_sc_hd__a221o_1 _0862_ (.A1(_0069_),
    .A2(_0206_),
    .B1(_0230_),
    .B2(_0375_),
    .C1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__xor2_1 _0863_ (.A(\game.v[4] ),
    .B(\game.paddle[4] ),
    .X(_0380_));
 sky130_fd_sc_hd__a221o_1 _0864_ (.A1(_0068_),
    .A2(_0203_),
    .B1(_0374_),
    .B2(_0104_),
    .C1(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__or4_1 _0865_ (.A(_0162_),
    .B(_0377_),
    .C(_0379_),
    .D(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__xor2_1 _0866_ (.A(_0088_),
    .B(\game.paddle[7] ),
    .X(_0383_));
 sky130_fd_sc_hd__a21oi_1 _0867_ (.A1(_0089_),
    .A2(_0243_),
    .B1(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__xnor2_1 _0868_ (.A(_0079_),
    .B(_0192_),
    .Y(_0385_));
 sky130_fd_sc_hd__or2_1 _0869_ (.A(_0089_),
    .B(_0243_),
    .X(_0386_));
 sky130_fd_sc_hd__and4b_1 _0870_ (.A_N(_0382_),
    .B(_0384_),
    .C(_0385_),
    .D(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__and3_1 _0871_ (.A(\game.inBallY ),
    .B(\game.inBallX ),
    .C(_0063_),
    .X(_0388_));
 sky130_fd_sc_hd__a21o_1 _0872_ (.A1(_0188_),
    .A2(\game.hit ),
    .B1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__and3b_1 _0873_ (.A_N(_0387_),
    .B(_0389_),
    .C(_0178_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _0874_ (.A(_0390_),
    .X(_0031_));
 sky130_fd_sc_hd__a211o_1 _0875_ (.A1(_0154_),
    .A2(_0155_),
    .B1(_0152_),
    .C1(_0153_),
    .X(_0391_));
 sky130_fd_sc_hd__xnor2_1 _0876_ (.A(_0060_),
    .B(\game.ballX[8] ),
    .Y(_0392_));
 sky130_fd_sc_hd__and3_1 _0877_ (.A(\game.ballX[3] ),
    .B(_0154_),
    .C(_0155_),
    .X(_0393_));
 sky130_fd_sc_hd__and2_1 _0878_ (.A(_0152_),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _0879_ (.A(\game.h[2] ),
    .B(\game.ballX[1] ),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _0880_ (.A(\game.h[2] ),
    .B(\game.ballX[1] ),
    .Y(_0396_));
 sky130_fd_sc_hd__nand2_1 _0881_ (.A(_0072_),
    .B(_0314_),
    .Y(_0397_));
 sky130_fd_sc_hd__or2_1 _0882_ (.A(_0072_),
    .B(_0314_),
    .X(_0398_));
 sky130_fd_sc_hd__a22o_1 _0883_ (.A1(_0395_),
    .A2(_0396_),
    .B1(_0397_),
    .B2(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__xor2_1 _0884_ (.A(_0073_),
    .B(\game.ballX[2] ),
    .X(_0400_));
 sky130_fd_sc_hd__xnor2_1 _0885_ (.A(_0061_),
    .B(\game.ballX[7] ),
    .Y(_0401_));
 sky130_fd_sc_hd__xnor2_1 _0886_ (.A(\game.h[4] ),
    .B(\game.ballX[3] ),
    .Y(_0402_));
 sky130_fd_sc_hd__xnor2_1 _0887_ (.A(\game.h[6] ),
    .B(_0155_),
    .Y(_0403_));
 sky130_fd_sc_hd__xnor2_1 _0888_ (.A(\game.h[7] ),
    .B(\game.ballX[6] ),
    .Y(_0404_));
 sky130_fd_sc_hd__and4_1 _0889_ (.A(_0401_),
    .B(_0402_),
    .C(_0403_),
    .D(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__xnor2_1 _0890_ (.A(_0099_),
    .B(_0154_),
    .Y(_0406_));
 sky130_fd_sc_hd__and4bb_1 _0891_ (.A_N(_0399_),
    .B_N(_0400_),
    .C(_0405_),
    .D(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__a31o_1 _0892_ (.A1(\game.inBallX ),
    .A2(_0153_),
    .A3(_0394_),
    .B1(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__xnor2_1 _0893_ (.A(_0394_),
    .B(_0401_),
    .Y(_0409_));
 sky130_fd_sc_hd__nor2_1 _0894_ (.A(\game.ballX[3] ),
    .B(_0154_),
    .Y(_0410_));
 sky130_fd_sc_hd__o21ai_1 _0895_ (.A1(\game.h[5] ),
    .A2(_0410_),
    .B1(_0403_),
    .Y(_0411_));
 sky130_fd_sc_hd__o31a_1 _0896_ (.A1(_0331_),
    .A2(_0344_),
    .A3(_0403_),
    .B1(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _0897_ (.A(_0331_),
    .B(_0344_),
    .Y(_0413_));
 sky130_fd_sc_hd__o21a_1 _0898_ (.A1(_0410_),
    .A2(_0413_),
    .B1(\game.h[5] ),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_1 _0899_ (.A(_0393_),
    .B(_0404_),
    .Y(_0415_));
 sky130_fd_sc_hd__or4_1 _0900_ (.A(_0399_),
    .B(_0402_),
    .C(_0414_),
    .D(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__a21oi_1 _0901_ (.A1(_0153_),
    .A2(_0394_),
    .B1(_0392_),
    .Y(_0417_));
 sky130_fd_sc_hd__a2111o_1 _0902_ (.A1(_0393_),
    .A2(_0404_),
    .B1(_0412_),
    .C1(_0416_),
    .D1(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__o31a_1 _0903_ (.A1(_0409_),
    .A2(_0400_),
    .A3(_0418_),
    .B1(\game.inBallX ),
    .X(_0419_));
 sky130_fd_sc_hd__a21oi_1 _0904_ (.A1(_0392_),
    .A2(_0408_),
    .B1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__a211oi_1 _0905_ (.A1(\game.ballX[8] ),
    .A2(_0391_),
    .B1(_0420_),
    .C1(_0267_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2_1 _0906_ (.A(\game.inBallY ),
    .B(_0081_),
    .Y(_0421_));
 sky130_fd_sc_hd__a21o_1 _0907_ (.A1(\game.inBallY ),
    .A2(_0085_),
    .B1(_0292_),
    .X(_0422_));
 sky130_fd_sc_hd__a21o_1 _0908_ (.A1(_0421_),
    .A2(_0422_),
    .B1(net23),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _0909_ (.A(\game.inBallX ),
    .B(_0083_),
    .Y(_0423_));
 sky130_fd_sc_hd__a211o_1 _0910_ (.A1(_0325_),
    .A2(_0423_),
    .B1(_0388_),
    .C1(_0267_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_2 _0911_ (.A(_0169_),
    .X(_0424_));
 sky130_fd_sc_hd__or2b_1 _0912_ (.A(_0089_),
    .B_N(_0144_),
    .X(_0425_));
 sky130_fd_sc_hd__or2b_1 _0913_ (.A(\game.ballY[5] ),
    .B_N(_0089_),
    .X(_0426_));
 sky130_fd_sc_hd__nand2_1 _0914_ (.A(_0090_),
    .B(_0289_),
    .Y(_0427_));
 sky130_fd_sc_hd__nand2_1 _0915_ (.A(_0375_),
    .B(\game.ballY[4] ),
    .Y(_0428_));
 sky130_fd_sc_hd__and4_1 _0916_ (.A(_0425_),
    .B(_0426_),
    .C(_0427_),
    .D(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_1 _0917_ (.A(_0066_),
    .B(_0255_),
    .Y(_0430_));
 sky130_fd_sc_hd__or2_1 _0918_ (.A(_0066_),
    .B(_0255_),
    .X(_0431_));
 sky130_fd_sc_hd__xor2_1 _0919_ (.A(_0095_),
    .B(\game.ballY[1] ),
    .X(_0432_));
 sky130_fd_sc_hd__a21oi_1 _0920_ (.A1(_0430_),
    .A2(_0431_),
    .B1(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__xor2_1 _0921_ (.A(_0104_),
    .B(\game.ballY[2] ),
    .X(_0434_));
 sky130_fd_sc_hd__xnor2_1 _0922_ (.A(_0127_),
    .B(_0149_),
    .Y(_0435_));
 sky130_fd_sc_hd__xnor2_1 _0923_ (.A(_0079_),
    .B(\game.ballY[7] ),
    .Y(_0436_));
 sky130_fd_sc_hd__xnor2_1 _0924_ (.A(_0088_),
    .B(\game.ballY[6] ),
    .Y(_0437_));
 sky130_fd_sc_hd__and4b_1 _0925_ (.A_N(_0434_),
    .B(_0435_),
    .C(_0436_),
    .D(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__a41o_1 _0926_ (.A1(_0424_),
    .A2(_0429_),
    .A3(_0433_),
    .A4(_0438_),
    .B1(\game.inBallY ),
    .X(_0439_));
 sky130_fd_sc_hd__nand3b_1 _0927_ (.A_N(_0427_),
    .B(_0426_),
    .C(_0425_),
    .Y(_0440_));
 sky130_fd_sc_hd__and3_1 _0928_ (.A(_0144_),
    .B(_0146_),
    .C(_0150_),
    .X(_0441_));
 sky130_fd_sc_hd__nand2_1 _0929_ (.A(_0147_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__a32o_1 _0930_ (.A1(_0149_),
    .A2(_0428_),
    .A3(_0440_),
    .B1(_0442_),
    .B2(_0080_),
    .X(_0443_));
 sky130_fd_sc_hd__a2bb2o_1 _0931_ (.A1_N(_0080_),
    .A2_N(_0442_),
    .B1(_0436_),
    .B2(_0441_),
    .X(_0444_));
 sky130_fd_sc_hd__a21o_1 _0932_ (.A1(_0144_),
    .A2(_0150_),
    .B1(_0437_),
    .X(_0445_));
 sky130_fd_sc_hd__inv_2 _0933_ (.A(\game.inBallY ),
    .Y(_0446_));
 sky130_fd_sc_hd__nor3_1 _0934_ (.A(_0446_),
    .B(_0434_),
    .C(_0435_),
    .Y(_0447_));
 sky130_fd_sc_hd__and4_1 _0935_ (.A(_0169_),
    .B(_0433_),
    .C(_0445_),
    .D(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__o211ai_1 _0936_ (.A1(_0437_),
    .A2(_0425_),
    .B1(_0426_),
    .C1(_0150_),
    .Y(_0449_));
 sky130_fd_sc_hd__o221a_1 _0937_ (.A1(_0441_),
    .A2(_0436_),
    .B1(_0429_),
    .B2(_0149_),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__or4bb_1 _0938_ (.A(_0443_),
    .B(_0444_),
    .C_N(_0448_),
    .D_N(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__and3_1 _0939_ (.A(_0175_),
    .B(_0439_),
    .C(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _0940_ (.A(_0452_),
    .X(_0035_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0941_ (.A(\game.h[0] ),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _0942_ (.A(_0058_),
    .B(_0169_),
    .Y(_0454_));
 sky130_fd_sc_hd__clkbuf_2 _0943_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__and2b_1 _0944_ (.A_N(_0453_),
    .B(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0945_ (.A(_0456_),
    .X(_0036_));
 sky130_fd_sc_hd__a21boi_1 _0946_ (.A1(_0076_),
    .A2(_0453_),
    .B1_N(_0454_),
    .Y(_0457_));
 sky130_fd_sc_hd__o21a_1 _0947_ (.A1(_0076_),
    .A2(_0453_),
    .B1(_0457_),
    .X(_0037_));
 sky130_fd_sc_hd__nand3_1 _0948_ (.A(_0076_),
    .B(_0453_),
    .C(_0074_),
    .Y(_0458_));
 sky130_fd_sc_hd__a21o_1 _0949_ (.A1(_0076_),
    .A2(_0453_),
    .B1(_0074_),
    .X(_0459_));
 sky130_fd_sc_hd__and3_1 _0950_ (.A(_0458_),
    .B(_0454_),
    .C(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(_0460_),
    .X(_0038_));
 sky130_fd_sc_hd__a31o_1 _0952_ (.A1(_0076_),
    .A2(_0453_),
    .A3(_0074_),
    .B1(_0073_),
    .X(_0461_));
 sky130_fd_sc_hd__and3b_1 _0953_ (.A_N(_0160_),
    .B(_0461_),
    .C(_0178_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _0954_ (.A(_0462_),
    .X(_0039_));
 sky130_fd_sc_hd__o21ai_1 _0955_ (.A1(_0077_),
    .A2(_0160_),
    .B1(_0245_),
    .Y(_0463_));
 sky130_fd_sc_hd__nor2_1 _0956_ (.A(_0161_),
    .B(_0463_),
    .Y(_0040_));
 sky130_fd_sc_hd__o21ai_1 _0957_ (.A1(_0099_),
    .A2(_0161_),
    .B1(_0455_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21oi_1 _0958_ (.A1(_0099_),
    .A2(_0161_),
    .B1(_0464_),
    .Y(_0041_));
 sky130_fd_sc_hd__and2_1 _0959_ (.A(_0100_),
    .B(_0160_),
    .X(_0465_));
 sky130_fd_sc_hd__a31o_1 _0960_ (.A1(_0099_),
    .A2(_0077_),
    .A3(_0160_),
    .B1(\game.h[6] ),
    .X(_0466_));
 sky130_fd_sc_hd__and3b_1 _0961_ (.A_N(_0465_),
    .B(_0454_),
    .C(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0962_ (.A(_0467_),
    .X(_0042_));
 sky130_fd_sc_hd__and3_1 _0963_ (.A(\game.h[7] ),
    .B(_0100_),
    .C(_0160_),
    .X(_0468_));
 sky130_fd_sc_hd__o21ai_1 _0964_ (.A1(\game.h[7] ),
    .A2(_0465_),
    .B1(_0455_),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_1 _0965_ (.A(_0468_),
    .B(_0469_),
    .Y(_0043_));
 sky130_fd_sc_hd__and2_1 _0966_ (.A(_0061_),
    .B(_0468_),
    .X(_0470_));
 sky130_fd_sc_hd__o21ai_1 _0967_ (.A1(_0061_),
    .A2(_0468_),
    .B1(_0455_),
    .Y(_0471_));
 sky130_fd_sc_hd__nor2_1 _0968_ (.A(_0470_),
    .B(_0471_),
    .Y(_0044_));
 sky130_fd_sc_hd__a21boi_1 _0969_ (.A1(_0060_),
    .A2(_0470_),
    .B1_N(_0454_),
    .Y(_0472_));
 sky130_fd_sc_hd__o21a_1 _0970_ (.A1(_0060_),
    .A2(_0470_),
    .B1(_0472_),
    .X(_0045_));
 sky130_fd_sc_hd__and3_1 _0971_ (.A(\game.paddle[6] ),
    .B(_0246_),
    .C(_0192_),
    .X(_0473_));
 sky130_fd_sc_hd__xnor2_1 _0972_ (.A(_0096_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _0973_ (.A(_0240_),
    .B(_0246_),
    .Y(_0475_));
 sky130_fd_sc_hd__xor2_1 _0974_ (.A(_0475_),
    .B(_0385_),
    .X(_0476_));
 sky130_fd_sc_hd__a21o_1 _0975_ (.A1(_0383_),
    .A2(_0386_),
    .B1(_0384_),
    .X(_0477_));
 sky130_fd_sc_hd__o41a_1 _0976_ (.A1(_0382_),
    .A2(_0474_),
    .A3(_0476_),
    .A4(_0477_),
    .B1(\game.inPaddle ),
    .X(_0478_));
 sky130_fd_sc_hd__o21a_1 _0977_ (.A1(_0387_),
    .A2(_0478_),
    .B1(_0176_),
    .X(_0046_));
 sky130_fd_sc_hd__nor2_1 _0978_ (.A(_0162_),
    .B(_0190_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0131_),
    .B(_0424_),
    .Y(_0480_));
 sky130_fd_sc_hd__o211a_1 _0980_ (.A1(_0131_),
    .A2(_0479_),
    .B1(_0480_),
    .C1(_0245_),
    .X(_0047_));
 sky130_fd_sc_hd__a31o_1 _0981_ (.A1(_0066_),
    .A2(_0131_),
    .A3(_0424_),
    .B1(_0059_),
    .X(_0481_));
 sky130_fd_sc_hd__a21oi_1 _0982_ (.A1(_0068_),
    .A2(_0480_),
    .B1(_0481_),
    .Y(_0048_));
 sky130_fd_sc_hd__and3_1 _0983_ (.A(\game.v[2] ),
    .B(_0065_),
    .C(\game.v[0] ),
    .X(_0482_));
 sky130_fd_sc_hd__a21oi_1 _0984_ (.A1(_0066_),
    .A2(_0131_),
    .B1(_0095_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_1 _0985_ (.A(_0482_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__a32o_1 _0986_ (.A1(_0245_),
    .A2(_0479_),
    .A3(_0484_),
    .B1(_0455_),
    .B2(_0095_),
    .X(_0049_));
 sky130_fd_sc_hd__nor2_1 _0987_ (.A(_0104_),
    .B(_0482_),
    .Y(_0485_));
 sky130_fd_sc_hd__and2_1 _0988_ (.A(\game.v[3] ),
    .B(_0482_),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_1 _0989_ (.A(_0485_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__a32o_1 _0990_ (.A1(_0245_),
    .A2(_0479_),
    .A3(_0487_),
    .B1(_0455_),
    .B2(_0104_),
    .X(_0050_));
 sky130_fd_sc_hd__and3_1 _0991_ (.A(_0127_),
    .B(_0169_),
    .C(_0486_),
    .X(_0488_));
 sky130_fd_sc_hd__a21o_1 _0992_ (.A1(_0424_),
    .A2(_0486_),
    .B1(_0127_),
    .X(_0489_));
 sky130_fd_sc_hd__and3b_1 _0993_ (.A_N(_0488_),
    .B(_0178_),
    .C(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(_0490_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _0995_ (.A(_0090_),
    .B(_0488_),
    .X(_0491_));
 sky130_fd_sc_hd__o21ai_1 _0996_ (.A1(_0090_),
    .A2(_0488_),
    .B1(_0200_),
    .Y(_0492_));
 sky130_fd_sc_hd__nor2_1 _0997_ (.A(_0491_),
    .B(_0492_),
    .Y(_0052_));
 sky130_fd_sc_hd__o21ai_1 _0998_ (.A1(_0159_),
    .A2(_0491_),
    .B1(_0200_),
    .Y(_0493_));
 sky130_fd_sc_hd__a21oi_1 _0999_ (.A1(_0159_),
    .A2(_0491_),
    .B1(_0493_),
    .Y(_0053_));
 sky130_fd_sc_hd__a31o_1 _1000_ (.A1(_0159_),
    .A2(_0090_),
    .A3(_0488_),
    .B1(_0088_),
    .X(_0494_));
 sky130_fd_sc_hd__nand3_1 _1001_ (.A(_0088_),
    .B(_0159_),
    .C(_0491_),
    .Y(_0495_));
 sky130_fd_sc_hd__and3_1 _1002_ (.A(_0175_),
    .B(_0494_),
    .C(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(_0496_),
    .X(_0054_));
 sky130_fd_sc_hd__a31o_1 _1004_ (.A1(_0088_),
    .A2(_0159_),
    .A3(_0491_),
    .B1(_0079_),
    .X(_0497_));
 sky130_fd_sc_hd__nand4_1 _1005_ (.A(_0127_),
    .B(_0091_),
    .C(_0424_),
    .D(_0486_),
    .Y(_0498_));
 sky130_fd_sc_hd__and3_1 _1006_ (.A(_0175_),
    .B(_0497_),
    .C(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(_0499_),
    .X(_0055_));
 sky130_fd_sc_hd__a31o_1 _1008_ (.A1(_0127_),
    .A2(_0091_),
    .A3(_0486_),
    .B1(_0165_),
    .X(_0500_));
 sky130_fd_sc_hd__and3_1 _1009_ (.A(_0080_),
    .B(_0424_),
    .C(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__a211oi_1 _1010_ (.A1(_0096_),
    .A2(_0498_),
    .B1(_0501_),
    .C1(_0267_),
    .Y(_0056_));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(net28),
    .D(_0000_),
    .Q(\game.offset[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(net37),
    .D(_0001_),
    .Q(\game.offset[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(net37),
    .D(_0002_),
    .Q(\game.offset[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(net38),
    .D(_0003_),
    .Q(\game.offset[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(net37),
    .D(_0004_),
    .Q(\game.offset[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(net33),
    .D(_0005_),
    .Q(\game.paddle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(net25),
    .D(_0006_),
    .Q(\game.paddle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(net31),
    .D(_0007_),
    .Q(\game.paddle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(net25),
    .D(_0008_),
    .Q(\game.paddle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(net26),
    .D(_0009_),
    .Q(\game.paddle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(net31),
    .D(_0010_),
    .Q(\game.paddle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(net33),
    .D(_0011_),
    .Q(\game.paddle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(net31),
    .D(_0012_),
    .Q(\game.paddle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(net31),
    .D(_0013_),
    .Q(\game.paddle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(net27),
    .D(_0014_),
    .Q(\game.ballY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(net28),
    .D(_0015_),
    .Q(\game.ballY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(net27),
    .D(_0016_),
    .Q(\game.ballY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(net27),
    .D(_0017_),
    .Q(\game.ballY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(net27),
    .D(_0018_),
    .Q(\game.ballY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(net29),
    .D(_0019_),
    .Q(\game.ballY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(net29),
    .D(_0020_),
    .Q(\game.ballY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(net29),
    .D(_0021_),
    .Q(\game.ballY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(net27),
    .D(_0022_),
    .Q(\game.ballX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(net28),
    .D(_0023_),
    .Q(\game.ballX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(net27),
    .D(_0024_),
    .Q(\game.ballX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(net25),
    .D(_0025_),
    .Q(\game.ballX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(net25),
    .D(_0026_),
    .Q(\game.ballX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(net25),
    .D(_0027_),
    .Q(\game.ballX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(net26),
    .D(_0028_),
    .Q(\game.ballX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(net26),
    .D(_0029_),
    .Q(\game.ballX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(net25),
    .D(_0030_),
    .Q(\game.ballX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(net35),
    .D(_0031_),
    .Q(\game.hit ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(net28),
    .D(_0032_),
    .Q(\game.inBallX ));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(net28),
    .D(_0033_),
    .Q(\game.ballDirY ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(net28),
    .D(_0034_),
    .Q(\game.ballDirX ));
 sky130_fd_sc_hd__dfxtp_2 _1046_ (.CLK(net35),
    .D(_0035_),
    .Q(\game.inBallY ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(net32),
    .D(_0036_),
    .Q(\game.h[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(net32),
    .D(_0037_),
    .Q(\game.h[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(net32),
    .D(_0038_),
    .Q(\game.h[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(net37),
    .D(_0039_),
    .Q(\game.h[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(net32),
    .D(_0040_),
    .Q(\game.h[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(net31),
    .D(_0041_),
    .Q(\game.h[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(net33),
    .D(_0042_),
    .Q(\game.h[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(net33),
    .D(_0043_),
    .Q(\game.h[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(net32),
    .D(_0044_),
    .Q(\game.h[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(net31),
    .D(_0045_),
    .Q(\game.h[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(net34),
    .D(_0046_),
    .Q(\game.inPaddle ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(net32),
    .D(_0047_),
    .Q(\game.v[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(net35),
    .D(_0048_),
    .Q(\game.v[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(net37),
    .D(_0049_),
    .Q(\game.v[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(net37),
    .D(_0050_),
    .Q(\game.v[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1062_ (.CLK(net35),
    .D(_0051_),
    .Q(\game.v[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(net35),
    .D(_0052_),
    .Q(\game.v[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(net36),
    .D(_0053_),
    .Q(\game.v[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(net36),
    .D(_0054_),
    .Q(\game.v[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(net36),
    .D(_0055_),
    .Q(\game.v[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(net35),
    .D(_0056_),
    .Q(\game.v[9] ));
 sky130_fd_sc_hd__conb_1 solo_squash_caravel_41 (.LO(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net10));
 sky130_fd_sc_hd__clkbuf_1 _1070_ (.A(net3),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 _1071_ (.A(net24),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 _1072_ (.A(net24),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 _1073_ (.A(net24),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 _1074_ (.A(net24),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 _1075_ (.A(net23),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 _1076_ (.A(net10),
    .X(net17));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(down_key_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ext_reset_n),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(gpio_ready),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(new_game_n),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(pause_n),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(up_key_n),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(wb_clk_i),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(wb_rst_i),
    .X(net8));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(blue));
 sky130_fd_sc_hd__buf_2 output10 (.A(net23),
    .X(debug_design_reset));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(debug_gpio_ready));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(design_oeb[0]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(design_oeb[1]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(design_oeb[2]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(design_oeb[3]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(design_oeb[4]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(design_oeb[5]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(green));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(hsync));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(red));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(speaker));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(vsync));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(net10),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(net30),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 fanout26 (.A(net30),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout27 (.A(net29),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout30 (.A(net39),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 fanout31 (.A(net34),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 fanout34 (.A(net39),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(net38),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 fanout36 (.A(net38),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout39 (.A(net7),
    .X(net39));
 sky130_fd_sc_hd__conb_1 solo_squash_caravel_40 (.LO(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net24));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
 assign debug_oeb[0] = net40;
 assign debug_oeb[1] = net41;
endmodule

